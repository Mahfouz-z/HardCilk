module stealNetworkDataUnit(
  input          clock,
  input          reset,
  input  [255:0] io_taskIn,
  output [255:0] io_taskOut,
  input          io_validIn,
  output         io_validOut,
  input          io_connSS_availableTask_ready,
  output         io_connSS_availableTask_valid,
  output [255:0] io_connSS_availableTask_bits,
  output         io_connSS_qOutTask_ready,
  input          io_connSS_qOutTask_valid,
  input  [255:0] io_connSS_qOutTask_bits,
  output         io_occupied
);
`ifdef RANDOMIZE_REG_INIT
  reg [255:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [255:0] taskReg; // @[stealNetworkDataUnit.scala 32:33]
  reg  validReg; // @[stealNetworkDataUnit.scala 33:33]
  wire  _T_2 = io_connSS_qOutTask_valid & ~io_validIn; // @[stealNetworkDataUnit.scala 50:41]
  wire  _GEN_2 = io_connSS_qOutTask_valid & ~io_validIn | io_validIn; // @[stealNetworkDataUnit.scala 50:56 51:32]
  assign io_taskOut = taskReg; // @[stealNetworkDataUnit.scala 63:25]
  assign io_validOut = validReg; // @[stealNetworkDataUnit.scala 64:25]
  assign io_connSS_availableTask_valid = io_connSS_availableTask_ready & io_validIn; // @[stealNetworkDataUnit.scala 45:40]
  assign io_connSS_availableTask_bits = io_connSS_availableTask_ready & io_validIn ? io_taskIn : 256'h0; // @[stealNetworkDataUnit.scala 42:35 45:54 49:37]
  assign io_connSS_qOutTask_ready = io_connSS_availableTask_ready & io_validIn ? 1'h0 : _T_2; // @[stealNetworkDataUnit.scala 41:30 45:54]
  assign io_occupied = validReg; // @[stealNetworkDataUnit.scala 65:25]
  always @(posedge clock) begin
    if (reset) begin // @[stealNetworkDataUnit.scala 32:33]
      taskReg <= 256'h0; // @[stealNetworkDataUnit.scala 32:33]
    end else if (io_connSS_availableTask_ready & io_validIn) begin // @[stealNetworkDataUnit.scala 45:54]
      taskReg <= 256'h0; // @[stealNetworkDataUnit.scala 47:37]
    end else if (io_connSS_qOutTask_valid & ~io_validIn) begin // @[stealNetworkDataUnit.scala 50:56]
      taskReg <= io_connSS_qOutTask_bits; // @[stealNetworkDataUnit.scala 52:32]
    end else if (io_validIn) begin // @[stealNetworkDataUnit.scala 54:27]
      taskReg <= io_taskIn; // @[stealNetworkDataUnit.scala 56:19]
    end else begin
      taskReg <= 256'h0; // @[stealNetworkDataUnit.scala 59:22]
    end
    if (reset) begin // @[stealNetworkDataUnit.scala 33:33]
      validReg <= 1'h0; // @[stealNetworkDataUnit.scala 33:33]
    end else if (io_connSS_availableTask_ready & io_validIn) begin // @[stealNetworkDataUnit.scala 45:54]
      validReg <= 1'h0; // @[stealNetworkDataUnit.scala 46:37]
    end else begin
      validReg <= _GEN_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {8{`RANDOM}};
  taskReg = _RAND_0[255:0];
  _RAND_1 = {1{`RANDOM}};
  validReg = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module stealNetworkCtrlUnit(
  input   clock,
  input   reset,
  input   io_reqTaskIn,
  output  io_reqTaskOut,
  output  io_connSS_serveStealReq_ready,
  input   io_connSS_serveStealReq_valid,
  output  io_connSS_stealReq_ready,
  input   io_connSS_stealReq_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  stealReqReg; // @[stealNetworkCtrlUnit.scala 20:28]
  wire  _GEN_0 = io_connSS_serveStealReq_valid ? 1'h0 : stealReqReg; // @[stealNetworkCtrlUnit.scala 24:44 25:19 27:19]
  assign io_reqTaskOut = io_connSS_stealReq_valid | _GEN_0; // @[stealNetworkCtrlUnit.scala 22:33 23:19]
  assign io_connSS_serveStealReq_ready = stealReqReg; // @[stealNetworkCtrlUnit.scala 31:33]
  assign io_connSS_stealReq_ready = ~stealReqReg; // @[stealNetworkCtrlUnit.scala 30:36]
  always @(posedge clock) begin
    if (reset) begin // @[stealNetworkCtrlUnit.scala 20:28]
      stealReqReg <= 1'h0; // @[stealNetworkCtrlUnit.scala 20:28]
    end else begin
      stealReqReg <= io_reqTaskIn; // @[stealNetworkCtrlUnit.scala 32:33]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stealReqReg = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module stealNetwork(
  input          clock,
  input          reset,
  output         io_connSS_0_ctrl_serveStealReq_ready,
  input          io_connSS_0_ctrl_serveStealReq_valid,
  input          io_connSS_0_data_availableTask_ready,
  output         io_connSS_0_data_availableTask_valid,
  output [255:0] io_connSS_0_data_availableTask_bits,
  output         io_connSS_0_data_qOutTask_ready,
  input          io_connSS_0_data_qOutTask_valid,
  input  [255:0] io_connSS_0_data_qOutTask_bits,
  output         io_connSS_1_ctrl_serveStealReq_ready,
  input          io_connSS_1_ctrl_serveStealReq_valid,
  output         io_connSS_1_data_qOutTask_ready,
  input          io_connSS_1_data_qOutTask_valid,
  input  [255:0] io_connSS_1_data_qOutTask_bits,
  output         io_connSS_2_ctrl_serveStealReq_ready,
  input          io_connSS_2_ctrl_serveStealReq_valid,
  output         io_connSS_2_data_qOutTask_ready,
  input          io_connSS_2_data_qOutTask_valid,
  input  [255:0] io_connSS_2_data_qOutTask_bits,
  output         io_connSS_3_ctrl_serveStealReq_ready,
  input          io_connSS_3_ctrl_serveStealReq_valid,
  output         io_connSS_3_ctrl_stealReq_ready,
  input          io_connSS_3_ctrl_stealReq_valid,
  input          io_connSS_3_data_availableTask_ready,
  output         io_connSS_3_data_availableTask_valid,
  output [255:0] io_connSS_3_data_availableTask_bits,
  output         io_connSS_3_data_qOutTask_ready,
  input          io_connSS_3_data_qOutTask_valid,
  input  [255:0] io_connSS_3_data_qOutTask_bits,
  output         io_connSS_4_ctrl_serveStealReq_ready,
  input          io_connSS_4_ctrl_serveStealReq_valid,
  output         io_connSS_4_ctrl_stealReq_ready,
  input          io_connSS_4_ctrl_stealReq_valid,
  input          io_connSS_4_data_availableTask_ready,
  output         io_connSS_4_data_availableTask_valid,
  output [255:0] io_connSS_4_data_availableTask_bits,
  output         io_connSS_4_data_qOutTask_ready,
  input          io_connSS_4_data_qOutTask_valid,
  input  [255:0] io_connSS_4_data_qOutTask_bits,
  output         io_connSS_5_ctrl_serveStealReq_ready,
  input          io_connSS_5_ctrl_serveStealReq_valid,
  output         io_connSS_5_ctrl_stealReq_ready,
  input          io_connSS_5_ctrl_stealReq_valid,
  input          io_connSS_5_data_availableTask_ready,
  output         io_connSS_5_data_availableTask_valid,
  output [255:0] io_connSS_5_data_availableTask_bits,
  output         io_connSS_5_data_qOutTask_ready,
  input          io_connSS_5_data_qOutTask_valid,
  input  [255:0] io_connSS_5_data_qOutTask_bits,
  output         io_connSS_6_ctrl_serveStealReq_ready,
  input          io_connSS_6_ctrl_serveStealReq_valid,
  output         io_connSS_6_ctrl_stealReq_ready,
  input          io_connSS_6_ctrl_stealReq_valid,
  input          io_connSS_6_data_availableTask_ready,
  output         io_connSS_6_data_availableTask_valid,
  output [255:0] io_connSS_6_data_availableTask_bits,
  output         io_connSS_6_data_qOutTask_ready,
  input          io_connSS_6_data_qOutTask_valid,
  input  [255:0] io_connSS_6_data_qOutTask_bits,
  output         io_connSS_7_ctrl_serveStealReq_ready,
  input          io_connSS_7_ctrl_serveStealReq_valid,
  output         io_connSS_7_ctrl_stealReq_ready,
  input          io_connSS_7_ctrl_stealReq_valid,
  input          io_connSS_7_data_availableTask_ready,
  output         io_connSS_7_data_availableTask_valid,
  output [255:0] io_connSS_7_data_availableTask_bits,
  output         io_connSS_7_data_qOutTask_ready,
  input          io_connSS_7_data_qOutTask_valid,
  input  [255:0] io_connSS_7_data_qOutTask_bits,
  output         io_connSS_8_ctrl_serveStealReq_ready,
  input          io_connSS_8_ctrl_serveStealReq_valid,
  output         io_connSS_8_ctrl_stealReq_ready,
  input          io_connSS_8_ctrl_stealReq_valid,
  input          io_connSS_8_data_availableTask_ready,
  output         io_connSS_8_data_availableTask_valid,
  output [255:0] io_connSS_8_data_availableTask_bits,
  output         io_connSS_8_data_qOutTask_ready,
  input          io_connSS_8_data_qOutTask_valid,
  input  [255:0] io_connSS_8_data_qOutTask_bits,
  output         io_connSS_9_ctrl_serveStealReq_ready,
  input          io_connSS_9_ctrl_serveStealReq_valid,
  output         io_connSS_9_ctrl_stealReq_ready,
  input          io_connSS_9_ctrl_stealReq_valid,
  input          io_connSS_9_data_availableTask_ready,
  output         io_connSS_9_data_availableTask_valid,
  output [255:0] io_connSS_9_data_availableTask_bits,
  output         io_connSS_9_data_qOutTask_ready,
  input          io_connSS_9_data_qOutTask_valid,
  input  [255:0] io_connSS_9_data_qOutTask_bits,
  output         io_connSS_10_ctrl_serveStealReq_ready,
  input          io_connSS_10_ctrl_serveStealReq_valid,
  output         io_connSS_10_ctrl_stealReq_ready,
  input          io_connSS_10_ctrl_stealReq_valid,
  input          io_connSS_10_data_availableTask_ready,
  output         io_connSS_10_data_availableTask_valid,
  output [255:0] io_connSS_10_data_availableTask_bits,
  output         io_connSS_10_data_qOutTask_ready,
  input          io_connSS_10_data_qOutTask_valid,
  input  [255:0] io_connSS_10_data_qOutTask_bits,
  output         io_connSS_11_ctrl_serveStealReq_ready,
  input          io_connSS_11_ctrl_serveStealReq_valid,
  output         io_connSS_11_ctrl_stealReq_ready,
  input          io_connSS_11_ctrl_stealReq_valid,
  input          io_connSS_11_data_availableTask_ready,
  output         io_connSS_11_data_availableTask_valid,
  output [255:0] io_connSS_11_data_availableTask_bits,
  output         io_connSS_11_data_qOutTask_ready,
  input          io_connSS_11_data_qOutTask_valid,
  input  [255:0] io_connSS_11_data_qOutTask_bits,
  output         io_connSS_12_ctrl_serveStealReq_ready,
  input          io_connSS_12_ctrl_serveStealReq_valid,
  output         io_connSS_12_ctrl_stealReq_ready,
  input          io_connSS_12_ctrl_stealReq_valid,
  input          io_connSS_12_data_availableTask_ready,
  output         io_connSS_12_data_availableTask_valid,
  output [255:0] io_connSS_12_data_availableTask_bits,
  output         io_connSS_12_data_qOutTask_ready,
  input          io_connSS_12_data_qOutTask_valid,
  input  [255:0] io_connSS_12_data_qOutTask_bits,
  output         io_connSS_13_ctrl_serveStealReq_ready,
  input          io_connSS_13_ctrl_serveStealReq_valid,
  output         io_connSS_13_ctrl_stealReq_ready,
  input          io_connSS_13_ctrl_stealReq_valid,
  input          io_connSS_13_data_availableTask_ready,
  output         io_connSS_13_data_availableTask_valid,
  output [255:0] io_connSS_13_data_availableTask_bits,
  output         io_connSS_13_data_qOutTask_ready,
  input          io_connSS_13_data_qOutTask_valid,
  input  [255:0] io_connSS_13_data_qOutTask_bits,
  output         io_connSS_14_ctrl_serveStealReq_ready,
  input          io_connSS_14_ctrl_serveStealReq_valid,
  output         io_connSS_14_ctrl_stealReq_ready,
  input          io_connSS_14_ctrl_stealReq_valid,
  input          io_connSS_14_data_availableTask_ready,
  output         io_connSS_14_data_availableTask_valid,
  output [255:0] io_connSS_14_data_availableTask_bits,
  output         io_connSS_14_data_qOutTask_ready,
  input          io_connSS_14_data_qOutTask_valid,
  input  [255:0] io_connSS_14_data_qOutTask_bits,
  output         io_connSS_15_ctrl_serveStealReq_ready,
  input          io_connSS_15_ctrl_serveStealReq_valid,
  output         io_connSS_15_ctrl_stealReq_ready,
  input          io_connSS_15_ctrl_stealReq_valid,
  input          io_connSS_15_data_availableTask_ready,
  output         io_connSS_15_data_availableTask_valid,
  output [255:0] io_connSS_15_data_availableTask_bits,
  output         io_connSS_15_data_qOutTask_ready,
  input          io_connSS_15_data_qOutTask_valid,
  input  [255:0] io_connSS_15_data_qOutTask_bits,
  output         io_connSS_16_ctrl_serveStealReq_ready,
  input          io_connSS_16_ctrl_serveStealReq_valid,
  output         io_connSS_16_ctrl_stealReq_ready,
  input          io_connSS_16_ctrl_stealReq_valid,
  input          io_connSS_16_data_availableTask_ready,
  output         io_connSS_16_data_availableTask_valid,
  output [255:0] io_connSS_16_data_availableTask_bits,
  output         io_connSS_16_data_qOutTask_ready,
  input          io_connSS_16_data_qOutTask_valid,
  input  [255:0] io_connSS_16_data_qOutTask_bits,
  output         io_connSS_17_ctrl_serveStealReq_ready,
  input          io_connSS_17_ctrl_serveStealReq_valid,
  output         io_connSS_17_ctrl_stealReq_ready,
  input          io_connSS_17_ctrl_stealReq_valid,
  input          io_connSS_17_data_availableTask_ready,
  output         io_connSS_17_data_availableTask_valid,
  output [255:0] io_connSS_17_data_availableTask_bits,
  output         io_connSS_17_data_qOutTask_ready,
  input          io_connSS_17_data_qOutTask_valid,
  input  [255:0] io_connSS_17_data_qOutTask_bits,
  output         io_connSS_18_ctrl_serveStealReq_ready,
  input          io_connSS_18_ctrl_serveStealReq_valid,
  output         io_connSS_18_ctrl_stealReq_ready,
  input          io_connSS_18_ctrl_stealReq_valid,
  input          io_connSS_18_data_availableTask_ready,
  output         io_connSS_18_data_availableTask_valid,
  output [255:0] io_connSS_18_data_availableTask_bits,
  output         io_connSS_18_data_qOutTask_ready,
  input          io_connSS_18_data_qOutTask_valid,
  input  [255:0] io_connSS_18_data_qOutTask_bits,
  output         io_connSS_19_ctrl_serveStealReq_ready,
  input          io_connSS_19_ctrl_serveStealReq_valid,
  output         io_connSS_19_ctrl_stealReq_ready,
  input          io_connSS_19_ctrl_stealReq_valid,
  input          io_connSS_19_data_availableTask_ready,
  output         io_connSS_19_data_availableTask_valid,
  output [255:0] io_connSS_19_data_availableTask_bits,
  output         io_connSS_19_data_qOutTask_ready,
  input          io_connSS_19_data_qOutTask_valid,
  input  [255:0] io_connSS_19_data_qOutTask_bits,
  output         io_connSS_20_ctrl_serveStealReq_ready,
  input          io_connSS_20_ctrl_serveStealReq_valid,
  output         io_connSS_20_ctrl_stealReq_ready,
  input          io_connSS_20_ctrl_stealReq_valid,
  input          io_connSS_20_data_availableTask_ready,
  output         io_connSS_20_data_availableTask_valid,
  output [255:0] io_connSS_20_data_availableTask_bits,
  output         io_connSS_20_data_qOutTask_ready,
  input          io_connSS_20_data_qOutTask_valid,
  input  [255:0] io_connSS_20_data_qOutTask_bits,
  output         io_connSS_21_ctrl_serveStealReq_ready,
  input          io_connSS_21_ctrl_serveStealReq_valid,
  output         io_connSS_21_ctrl_stealReq_ready,
  input          io_connSS_21_ctrl_stealReq_valid,
  input          io_connSS_21_data_availableTask_ready,
  output         io_connSS_21_data_availableTask_valid,
  output [255:0] io_connSS_21_data_availableTask_bits,
  output         io_connSS_21_data_qOutTask_ready,
  input          io_connSS_21_data_qOutTask_valid,
  input  [255:0] io_connSS_21_data_qOutTask_bits,
  output         io_connSS_22_ctrl_serveStealReq_ready,
  input          io_connSS_22_ctrl_serveStealReq_valid,
  output         io_connSS_22_ctrl_stealReq_ready,
  input          io_connSS_22_ctrl_stealReq_valid,
  input          io_connSS_22_data_availableTask_ready,
  output         io_connSS_22_data_availableTask_valid,
  output [255:0] io_connSS_22_data_availableTask_bits,
  output         io_connSS_22_data_qOutTask_ready,
  input          io_connSS_22_data_qOutTask_valid,
  input  [255:0] io_connSS_22_data_qOutTask_bits,
  output         io_connSS_23_ctrl_serveStealReq_ready,
  input          io_connSS_23_ctrl_serveStealReq_valid,
  output         io_connSS_23_ctrl_stealReq_ready,
  input          io_connSS_23_ctrl_stealReq_valid,
  input          io_connSS_23_data_availableTask_ready,
  output         io_connSS_23_data_availableTask_valid,
  output [255:0] io_connSS_23_data_availableTask_bits,
  output         io_connSS_23_data_qOutTask_ready,
  input          io_connSS_23_data_qOutTask_valid,
  input  [255:0] io_connSS_23_data_qOutTask_bits,
  output         io_connSS_24_ctrl_serveStealReq_ready,
  input          io_connSS_24_ctrl_serveStealReq_valid,
  output         io_connSS_24_ctrl_stealReq_ready,
  input          io_connSS_24_ctrl_stealReq_valid,
  input          io_connSS_24_data_availableTask_ready,
  output         io_connSS_24_data_availableTask_valid,
  output [255:0] io_connSS_24_data_availableTask_bits,
  output         io_connSS_24_data_qOutTask_ready,
  input          io_connSS_24_data_qOutTask_valid,
  input  [255:0] io_connSS_24_data_qOutTask_bits,
  output         io_connSS_25_ctrl_serveStealReq_ready,
  input          io_connSS_25_ctrl_serveStealReq_valid,
  output         io_connSS_25_ctrl_stealReq_ready,
  input          io_connSS_25_ctrl_stealReq_valid,
  input          io_connSS_25_data_availableTask_ready,
  output         io_connSS_25_data_availableTask_valid,
  output [255:0] io_connSS_25_data_availableTask_bits,
  output         io_connSS_25_data_qOutTask_ready,
  input          io_connSS_25_data_qOutTask_valid,
  input  [255:0] io_connSS_25_data_qOutTask_bits,
  output         io_connSS_26_ctrl_serveStealReq_ready,
  input          io_connSS_26_ctrl_serveStealReq_valid,
  output         io_connSS_26_ctrl_stealReq_ready,
  input          io_connSS_26_ctrl_stealReq_valid,
  input          io_connSS_26_data_availableTask_ready,
  output         io_connSS_26_data_availableTask_valid,
  output [255:0] io_connSS_26_data_availableTask_bits,
  output         io_connSS_26_data_qOutTask_ready,
  input          io_connSS_26_data_qOutTask_valid,
  input  [255:0] io_connSS_26_data_qOutTask_bits,
  output         io_connSS_27_ctrl_serveStealReq_ready,
  input          io_connSS_27_ctrl_serveStealReq_valid,
  output         io_connSS_27_ctrl_stealReq_ready,
  input          io_connSS_27_ctrl_stealReq_valid,
  input          io_connSS_27_data_availableTask_ready,
  output         io_connSS_27_data_availableTask_valid,
  output [255:0] io_connSS_27_data_availableTask_bits,
  output         io_connSS_27_data_qOutTask_ready,
  input          io_connSS_27_data_qOutTask_valid,
  input  [255:0] io_connSS_27_data_qOutTask_bits,
  output         io_connSS_28_ctrl_serveStealReq_ready,
  input          io_connSS_28_ctrl_serveStealReq_valid,
  output         io_connSS_28_ctrl_stealReq_ready,
  input          io_connSS_28_ctrl_stealReq_valid,
  input          io_connSS_28_data_availableTask_ready,
  output         io_connSS_28_data_availableTask_valid,
  output [255:0] io_connSS_28_data_availableTask_bits,
  output         io_connSS_28_data_qOutTask_ready,
  input          io_connSS_28_data_qOutTask_valid,
  input  [255:0] io_connSS_28_data_qOutTask_bits,
  output         io_connSS_29_ctrl_serveStealReq_ready,
  input          io_connSS_29_ctrl_serveStealReq_valid,
  output         io_connSS_29_ctrl_stealReq_ready,
  input          io_connSS_29_ctrl_stealReq_valid,
  input          io_connSS_29_data_availableTask_ready,
  output         io_connSS_29_data_availableTask_valid,
  output [255:0] io_connSS_29_data_availableTask_bits,
  output         io_connSS_29_data_qOutTask_ready,
  input          io_connSS_29_data_qOutTask_valid,
  input  [255:0] io_connSS_29_data_qOutTask_bits,
  output         io_connSS_30_ctrl_serveStealReq_ready,
  input          io_connSS_30_ctrl_serveStealReq_valid,
  output         io_connSS_30_ctrl_stealReq_ready,
  input          io_connSS_30_ctrl_stealReq_valid,
  input          io_connSS_30_data_availableTask_ready,
  output         io_connSS_30_data_availableTask_valid,
  output [255:0] io_connSS_30_data_availableTask_bits,
  output         io_connSS_30_data_qOutTask_ready,
  input          io_connSS_30_data_qOutTask_valid,
  input  [255:0] io_connSS_30_data_qOutTask_bits,
  output         io_connSS_31_ctrl_serveStealReq_ready,
  input          io_connSS_31_ctrl_serveStealReq_valid,
  output         io_connSS_31_ctrl_stealReq_ready,
  input          io_connSS_31_ctrl_stealReq_valid,
  input          io_connSS_31_data_availableTask_ready,
  output         io_connSS_31_data_availableTask_valid,
  output [255:0] io_connSS_31_data_availableTask_bits,
  output         io_connSS_31_data_qOutTask_ready,
  input          io_connSS_31_data_qOutTask_valid,
  input  [255:0] io_connSS_31_data_qOutTask_bits,
  output         io_connSS_32_ctrl_serveStealReq_ready,
  input          io_connSS_32_ctrl_serveStealReq_valid,
  output         io_connSS_32_ctrl_stealReq_ready,
  input          io_connSS_32_ctrl_stealReq_valid,
  input          io_connSS_32_data_availableTask_ready,
  output         io_connSS_32_data_availableTask_valid,
  output [255:0] io_connSS_32_data_availableTask_bits,
  output         io_connSS_32_data_qOutTask_ready,
  input          io_connSS_32_data_qOutTask_valid,
  input  [255:0] io_connSS_32_data_qOutTask_bits,
  output         io_connSS_33_ctrl_serveStealReq_ready,
  input          io_connSS_33_ctrl_serveStealReq_valid,
  output         io_connSS_33_ctrl_stealReq_ready,
  input          io_connSS_33_ctrl_stealReq_valid,
  input          io_connSS_33_data_availableTask_ready,
  output         io_connSS_33_data_availableTask_valid,
  output [255:0] io_connSS_33_data_availableTask_bits,
  output         io_connSS_33_data_qOutTask_ready,
  input          io_connSS_33_data_qOutTask_valid,
  input  [255:0] io_connSS_33_data_qOutTask_bits,
  output         io_connSS_34_ctrl_serveStealReq_ready,
  input          io_connSS_34_ctrl_serveStealReq_valid,
  output         io_connSS_34_ctrl_stealReq_ready,
  input          io_connSS_34_ctrl_stealReq_valid,
  input          io_connSS_34_data_availableTask_ready,
  output         io_connSS_34_data_availableTask_valid,
  output [255:0] io_connSS_34_data_availableTask_bits,
  output         io_connSS_34_data_qOutTask_ready,
  input          io_connSS_34_data_qOutTask_valid,
  input  [255:0] io_connSS_34_data_qOutTask_bits,
  output         io_connSS_35_ctrl_serveStealReq_ready,
  input          io_connSS_35_ctrl_serveStealReq_valid,
  output         io_connSS_35_ctrl_stealReq_ready,
  input          io_connSS_35_ctrl_stealReq_valid,
  input          io_connSS_35_data_availableTask_ready,
  output         io_connSS_35_data_availableTask_valid,
  output [255:0] io_connSS_35_data_availableTask_bits,
  output         io_connSS_35_data_qOutTask_ready,
  input          io_connSS_35_data_qOutTask_valid,
  input  [255:0] io_connSS_35_data_qOutTask_bits,
  output         io_connSS_36_ctrl_serveStealReq_ready,
  input          io_connSS_36_ctrl_serveStealReq_valid,
  output         io_connSS_36_ctrl_stealReq_ready,
  input          io_connSS_36_ctrl_stealReq_valid,
  input          io_connSS_36_data_availableTask_ready,
  output         io_connSS_36_data_availableTask_valid,
  output [255:0] io_connSS_36_data_availableTask_bits,
  output         io_connSS_36_data_qOutTask_ready,
  input          io_connSS_36_data_qOutTask_valid,
  input  [255:0] io_connSS_36_data_qOutTask_bits,
  output         io_connSS_37_ctrl_serveStealReq_ready,
  input          io_connSS_37_ctrl_serveStealReq_valid,
  output         io_connSS_37_ctrl_stealReq_ready,
  input          io_connSS_37_ctrl_stealReq_valid,
  input          io_connSS_37_data_availableTask_ready,
  output         io_connSS_37_data_availableTask_valid,
  output [255:0] io_connSS_37_data_availableTask_bits,
  output         io_connSS_37_data_qOutTask_ready,
  input          io_connSS_37_data_qOutTask_valid,
  input  [255:0] io_connSS_37_data_qOutTask_bits,
  output         io_connSS_38_ctrl_serveStealReq_ready,
  input          io_connSS_38_ctrl_serveStealReq_valid,
  output         io_connSS_38_ctrl_stealReq_ready,
  input          io_connSS_38_ctrl_stealReq_valid,
  input          io_connSS_38_data_availableTask_ready,
  output         io_connSS_38_data_availableTask_valid,
  output [255:0] io_connSS_38_data_availableTask_bits,
  output         io_connSS_38_data_qOutTask_ready,
  input          io_connSS_38_data_qOutTask_valid,
  input  [255:0] io_connSS_38_data_qOutTask_bits,
  output         io_connSS_39_ctrl_serveStealReq_ready,
  input          io_connSS_39_ctrl_serveStealReq_valid,
  output         io_connSS_39_ctrl_stealReq_ready,
  input          io_connSS_39_ctrl_stealReq_valid,
  input          io_connSS_39_data_availableTask_ready,
  output         io_connSS_39_data_availableTask_valid,
  output [255:0] io_connSS_39_data_availableTask_bits,
  output         io_connSS_39_data_qOutTask_ready,
  input          io_connSS_39_data_qOutTask_valid,
  input  [255:0] io_connSS_39_data_qOutTask_bits,
  output         io_connSS_40_ctrl_serveStealReq_ready,
  input          io_connSS_40_ctrl_serveStealReq_valid,
  output         io_connSS_40_ctrl_stealReq_ready,
  input          io_connSS_40_ctrl_stealReq_valid,
  input          io_connSS_40_data_availableTask_ready,
  output         io_connSS_40_data_availableTask_valid,
  output [255:0] io_connSS_40_data_availableTask_bits,
  output         io_connSS_40_data_qOutTask_ready,
  input          io_connSS_40_data_qOutTask_valid,
  input  [255:0] io_connSS_40_data_qOutTask_bits,
  output         io_connSS_41_ctrl_serveStealReq_ready,
  input          io_connSS_41_ctrl_serveStealReq_valid,
  output         io_connSS_41_ctrl_stealReq_ready,
  input          io_connSS_41_ctrl_stealReq_valid,
  input          io_connSS_41_data_availableTask_ready,
  output         io_connSS_41_data_availableTask_valid,
  output [255:0] io_connSS_41_data_availableTask_bits,
  output         io_connSS_41_data_qOutTask_ready,
  input          io_connSS_41_data_qOutTask_valid,
  input  [255:0] io_connSS_41_data_qOutTask_bits,
  output         io_connSS_42_ctrl_serveStealReq_ready,
  input          io_connSS_42_ctrl_serveStealReq_valid,
  output         io_connSS_42_ctrl_stealReq_ready,
  input          io_connSS_42_ctrl_stealReq_valid,
  input          io_connSS_42_data_availableTask_ready,
  output         io_connSS_42_data_availableTask_valid,
  output [255:0] io_connSS_42_data_availableTask_bits,
  output         io_connSS_42_data_qOutTask_ready,
  input          io_connSS_42_data_qOutTask_valid,
  input  [255:0] io_connSS_42_data_qOutTask_bits,
  output         io_connSS_43_ctrl_serveStealReq_ready,
  input          io_connSS_43_ctrl_serveStealReq_valid,
  output         io_connSS_43_ctrl_stealReq_ready,
  input          io_connSS_43_ctrl_stealReq_valid,
  input          io_connSS_43_data_availableTask_ready,
  output         io_connSS_43_data_availableTask_valid,
  output [255:0] io_connSS_43_data_availableTask_bits,
  output         io_connSS_43_data_qOutTask_ready,
  input          io_connSS_43_data_qOutTask_valid,
  input  [255:0] io_connSS_43_data_qOutTask_bits,
  output         io_connSS_44_ctrl_serveStealReq_ready,
  input          io_connSS_44_ctrl_serveStealReq_valid,
  output         io_connSS_44_ctrl_stealReq_ready,
  input          io_connSS_44_ctrl_stealReq_valid,
  input          io_connSS_44_data_availableTask_ready,
  output         io_connSS_44_data_availableTask_valid,
  output [255:0] io_connSS_44_data_availableTask_bits,
  output         io_connSS_44_data_qOutTask_ready,
  input          io_connSS_44_data_qOutTask_valid,
  input  [255:0] io_connSS_44_data_qOutTask_bits,
  output         io_connSS_45_ctrl_serveStealReq_ready,
  input          io_connSS_45_ctrl_serveStealReq_valid,
  output         io_connSS_45_ctrl_stealReq_ready,
  input          io_connSS_45_ctrl_stealReq_valid,
  input          io_connSS_45_data_availableTask_ready,
  output         io_connSS_45_data_availableTask_valid,
  output [255:0] io_connSS_45_data_availableTask_bits,
  output         io_connSS_45_data_qOutTask_ready,
  input          io_connSS_45_data_qOutTask_valid,
  input  [255:0] io_connSS_45_data_qOutTask_bits,
  output         io_connSS_46_ctrl_serveStealReq_ready,
  input          io_connSS_46_ctrl_serveStealReq_valid,
  output         io_connSS_46_ctrl_stealReq_ready,
  input          io_connSS_46_ctrl_stealReq_valid,
  input          io_connSS_46_data_availableTask_ready,
  output         io_connSS_46_data_availableTask_valid,
  output [255:0] io_connSS_46_data_availableTask_bits,
  output         io_connSS_46_data_qOutTask_ready,
  input          io_connSS_46_data_qOutTask_valid,
  input  [255:0] io_connSS_46_data_qOutTask_bits,
  output         io_connSS_47_ctrl_serveStealReq_ready,
  input          io_connSS_47_ctrl_serveStealReq_valid,
  output         io_connSS_47_ctrl_stealReq_ready,
  input          io_connSS_47_ctrl_stealReq_valid,
  input          io_connSS_47_data_availableTask_ready,
  output         io_connSS_47_data_availableTask_valid,
  output [255:0] io_connSS_47_data_availableTask_bits,
  output         io_connSS_47_data_qOutTask_ready,
  input          io_connSS_47_data_qOutTask_valid,
  input  [255:0] io_connSS_47_data_qOutTask_bits,
  output         io_connSS_48_ctrl_serveStealReq_ready,
  input          io_connSS_48_ctrl_serveStealReq_valid,
  output         io_connSS_48_ctrl_stealReq_ready,
  input          io_connSS_48_ctrl_stealReq_valid,
  input          io_connSS_48_data_availableTask_ready,
  output         io_connSS_48_data_availableTask_valid,
  output [255:0] io_connSS_48_data_availableTask_bits,
  output         io_connSS_48_data_qOutTask_ready,
  input          io_connSS_48_data_qOutTask_valid,
  input  [255:0] io_connSS_48_data_qOutTask_bits,
  output         io_connSS_49_ctrl_serveStealReq_ready,
  input          io_connSS_49_ctrl_serveStealReq_valid,
  output         io_connSS_49_ctrl_stealReq_ready,
  input          io_connSS_49_ctrl_stealReq_valid,
  input          io_connSS_49_data_availableTask_ready,
  output         io_connSS_49_data_availableTask_valid,
  output [255:0] io_connSS_49_data_availableTask_bits,
  output         io_connSS_49_data_qOutTask_ready,
  input          io_connSS_49_data_qOutTask_valid,
  input  [255:0] io_connSS_49_data_qOutTask_bits,
  output         io_connSS_50_ctrl_serveStealReq_ready,
  input          io_connSS_50_ctrl_serveStealReq_valid,
  output         io_connSS_50_ctrl_stealReq_ready,
  input          io_connSS_50_ctrl_stealReq_valid,
  input          io_connSS_50_data_availableTask_ready,
  output         io_connSS_50_data_availableTask_valid,
  output [255:0] io_connSS_50_data_availableTask_bits,
  output         io_connSS_50_data_qOutTask_ready,
  input          io_connSS_50_data_qOutTask_valid,
  input  [255:0] io_connSS_50_data_qOutTask_bits,
  output         io_connSS_51_ctrl_serveStealReq_ready,
  input          io_connSS_51_ctrl_serveStealReq_valid,
  output         io_connSS_51_ctrl_stealReq_ready,
  input          io_connSS_51_ctrl_stealReq_valid,
  input          io_connSS_51_data_availableTask_ready,
  output         io_connSS_51_data_availableTask_valid,
  output [255:0] io_connSS_51_data_availableTask_bits,
  output         io_connSS_51_data_qOutTask_ready,
  input          io_connSS_51_data_qOutTask_valid,
  input  [255:0] io_connSS_51_data_qOutTask_bits,
  output         io_connSS_52_ctrl_serveStealReq_ready,
  input          io_connSS_52_ctrl_serveStealReq_valid,
  output         io_connSS_52_ctrl_stealReq_ready,
  input          io_connSS_52_ctrl_stealReq_valid,
  input          io_connSS_52_data_availableTask_ready,
  output         io_connSS_52_data_availableTask_valid,
  output [255:0] io_connSS_52_data_availableTask_bits,
  output         io_connSS_52_data_qOutTask_ready,
  input          io_connSS_52_data_qOutTask_valid,
  input  [255:0] io_connSS_52_data_qOutTask_bits,
  output         io_connSS_53_ctrl_serveStealReq_ready,
  input          io_connSS_53_ctrl_serveStealReq_valid,
  output         io_connSS_53_ctrl_stealReq_ready,
  input          io_connSS_53_ctrl_stealReq_valid,
  input          io_connSS_53_data_availableTask_ready,
  output         io_connSS_53_data_availableTask_valid,
  output [255:0] io_connSS_53_data_availableTask_bits,
  output         io_connSS_53_data_qOutTask_ready,
  input          io_connSS_53_data_qOutTask_valid,
  input  [255:0] io_connSS_53_data_qOutTask_bits,
  output         io_connSS_54_ctrl_serveStealReq_ready,
  input          io_connSS_54_ctrl_serveStealReq_valid,
  output         io_connSS_54_ctrl_stealReq_ready,
  input          io_connSS_54_ctrl_stealReq_valid,
  input          io_connSS_54_data_availableTask_ready,
  output         io_connSS_54_data_availableTask_valid,
  output [255:0] io_connSS_54_data_availableTask_bits,
  output         io_connSS_54_data_qOutTask_ready,
  input          io_connSS_54_data_qOutTask_valid,
  input  [255:0] io_connSS_54_data_qOutTask_bits,
  output         io_connSS_55_ctrl_serveStealReq_ready,
  input          io_connSS_55_ctrl_serveStealReq_valid,
  output         io_connSS_55_ctrl_stealReq_ready,
  input          io_connSS_55_ctrl_stealReq_valid,
  input          io_connSS_55_data_availableTask_ready,
  output         io_connSS_55_data_availableTask_valid,
  output [255:0] io_connSS_55_data_availableTask_bits,
  output         io_connSS_55_data_qOutTask_ready,
  input          io_connSS_55_data_qOutTask_valid,
  input  [255:0] io_connSS_55_data_qOutTask_bits,
  output         io_connSS_56_ctrl_serveStealReq_ready,
  input          io_connSS_56_ctrl_serveStealReq_valid,
  output         io_connSS_56_ctrl_stealReq_ready,
  input          io_connSS_56_ctrl_stealReq_valid,
  input          io_connSS_56_data_availableTask_ready,
  output         io_connSS_56_data_availableTask_valid,
  output [255:0] io_connSS_56_data_availableTask_bits,
  output         io_connSS_56_data_qOutTask_ready,
  input          io_connSS_56_data_qOutTask_valid,
  input  [255:0] io_connSS_56_data_qOutTask_bits,
  output         io_connSS_57_ctrl_serveStealReq_ready,
  input          io_connSS_57_ctrl_serveStealReq_valid,
  output         io_connSS_57_ctrl_stealReq_ready,
  input          io_connSS_57_ctrl_stealReq_valid,
  input          io_connSS_57_data_availableTask_ready,
  output         io_connSS_57_data_availableTask_valid,
  output [255:0] io_connSS_57_data_availableTask_bits,
  output         io_connSS_57_data_qOutTask_ready,
  input          io_connSS_57_data_qOutTask_valid,
  input  [255:0] io_connSS_57_data_qOutTask_bits,
  output         io_connSS_58_ctrl_serveStealReq_ready,
  input          io_connSS_58_ctrl_serveStealReq_valid,
  output         io_connSS_58_ctrl_stealReq_ready,
  input          io_connSS_58_ctrl_stealReq_valid,
  input          io_connSS_58_data_availableTask_ready,
  output         io_connSS_58_data_availableTask_valid,
  output [255:0] io_connSS_58_data_availableTask_bits,
  output         io_connSS_58_data_qOutTask_ready,
  input          io_connSS_58_data_qOutTask_valid,
  input  [255:0] io_connSS_58_data_qOutTask_bits,
  output         io_connSS_59_ctrl_serveStealReq_ready,
  input          io_connSS_59_ctrl_serveStealReq_valid,
  output         io_connSS_59_ctrl_stealReq_ready,
  input          io_connSS_59_ctrl_stealReq_valid,
  input          io_connSS_59_data_availableTask_ready,
  output         io_connSS_59_data_availableTask_valid,
  output [255:0] io_connSS_59_data_availableTask_bits,
  output         io_connSS_59_data_qOutTask_ready,
  input          io_connSS_59_data_qOutTask_valid,
  input  [255:0] io_connSS_59_data_qOutTask_bits,
  output         io_connSS_60_ctrl_serveStealReq_ready,
  input          io_connSS_60_ctrl_serveStealReq_valid,
  output         io_connSS_60_ctrl_stealReq_ready,
  input          io_connSS_60_ctrl_stealReq_valid,
  input          io_connSS_60_data_availableTask_ready,
  output         io_connSS_60_data_availableTask_valid,
  output [255:0] io_connSS_60_data_availableTask_bits,
  output         io_connSS_60_data_qOutTask_ready,
  input          io_connSS_60_data_qOutTask_valid,
  input  [255:0] io_connSS_60_data_qOutTask_bits,
  output         io_connSS_61_ctrl_serveStealReq_ready,
  input          io_connSS_61_ctrl_serveStealReq_valid,
  output         io_connSS_61_ctrl_stealReq_ready,
  input          io_connSS_61_ctrl_stealReq_valid,
  input          io_connSS_61_data_availableTask_ready,
  output         io_connSS_61_data_availableTask_valid,
  output [255:0] io_connSS_61_data_availableTask_bits,
  output         io_connSS_61_data_qOutTask_ready,
  input          io_connSS_61_data_qOutTask_valid,
  input  [255:0] io_connSS_61_data_qOutTask_bits,
  output         io_connSS_62_ctrl_serveStealReq_ready,
  input          io_connSS_62_ctrl_serveStealReq_valid,
  output         io_connSS_62_ctrl_stealReq_ready,
  input          io_connSS_62_ctrl_stealReq_valid,
  input          io_connSS_62_data_availableTask_ready,
  output         io_connSS_62_data_availableTask_valid,
  output [255:0] io_connSS_62_data_availableTask_bits,
  output         io_connSS_62_data_qOutTask_ready,
  input          io_connSS_62_data_qOutTask_valid,
  input  [255:0] io_connSS_62_data_qOutTask_bits,
  output         io_connSS_63_ctrl_serveStealReq_ready,
  input          io_connSS_63_ctrl_serveStealReq_valid,
  output         io_connSS_63_ctrl_stealReq_ready,
  input          io_connSS_63_ctrl_stealReq_valid,
  input          io_connSS_63_data_availableTask_ready,
  output         io_connSS_63_data_availableTask_valid,
  output [255:0] io_connSS_63_data_availableTask_bits,
  output         io_connSS_63_data_qOutTask_ready,
  input          io_connSS_63_data_qOutTask_valid,
  input  [255:0] io_connSS_63_data_qOutTask_bits,
  output         io_connSS_64_ctrl_serveStealReq_ready,
  input          io_connSS_64_ctrl_serveStealReq_valid,
  output         io_connSS_64_ctrl_stealReq_ready,
  input          io_connSS_64_ctrl_stealReq_valid,
  input          io_connSS_64_data_availableTask_ready,
  output         io_connSS_64_data_availableTask_valid,
  output [255:0] io_connSS_64_data_availableTask_bits,
  output         io_connSS_64_data_qOutTask_ready,
  input          io_connSS_64_data_qOutTask_valid,
  input  [255:0] io_connSS_64_data_qOutTask_bits,
  output         io_connSS_65_ctrl_serveStealReq_ready,
  input          io_connSS_65_ctrl_serveStealReq_valid,
  output         io_connSS_65_ctrl_stealReq_ready,
  input          io_connSS_65_ctrl_stealReq_valid,
  input          io_connSS_65_data_availableTask_ready,
  output         io_connSS_65_data_availableTask_valid,
  output [255:0] io_connSS_65_data_availableTask_bits,
  output         io_connSS_65_data_qOutTask_ready,
  input          io_connSS_65_data_qOutTask_valid,
  input  [255:0] io_connSS_65_data_qOutTask_bits,
  output         io_connSS_66_ctrl_serveStealReq_ready,
  input          io_connSS_66_ctrl_serveStealReq_valid,
  output         io_connSS_66_ctrl_stealReq_ready,
  input          io_connSS_66_ctrl_stealReq_valid,
  input          io_connSS_66_data_availableTask_ready,
  output         io_connSS_66_data_availableTask_valid,
  output [255:0] io_connSS_66_data_availableTask_bits,
  output         io_connSS_66_data_qOutTask_ready,
  input          io_connSS_66_data_qOutTask_valid,
  input  [255:0] io_connSS_66_data_qOutTask_bits,
  output         io_ntwDataUnitOccupancyVSS_0
);
  wire  dataUnits_0_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_0_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_0_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_0_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_0_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_0_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_0_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_0_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_0_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_0_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_0_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_0_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_0_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_1_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_1_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_1_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_1_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_1_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_1_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_1_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_1_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_1_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_1_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_1_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_1_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_1_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_2_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_2_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_2_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_2_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_2_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_2_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_2_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_2_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_2_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_2_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_2_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_2_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_2_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_3_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_3_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_3_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_3_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_3_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_3_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_3_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_3_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_3_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_3_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_3_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_3_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_3_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_4_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_4_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_4_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_4_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_4_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_4_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_4_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_4_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_4_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_4_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_4_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_4_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_4_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_5_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_5_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_5_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_5_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_5_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_5_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_5_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_5_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_5_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_5_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_5_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_5_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_5_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_6_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_6_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_6_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_6_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_6_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_6_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_6_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_6_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_6_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_6_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_6_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_6_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_6_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_7_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_7_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_7_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_7_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_7_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_7_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_7_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_7_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_7_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_7_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_7_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_7_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_7_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_8_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_8_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_8_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_8_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_8_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_8_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_8_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_8_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_8_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_8_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_8_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_8_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_8_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_9_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_9_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_9_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_9_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_9_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_9_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_9_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_9_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_9_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_9_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_9_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_9_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_9_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_10_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_10_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_10_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_10_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_10_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_10_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_10_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_10_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_10_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_10_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_10_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_10_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_10_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_11_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_11_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_11_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_11_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_11_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_11_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_11_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_11_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_11_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_11_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_11_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_11_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_11_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_12_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_12_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_12_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_12_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_12_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_12_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_12_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_12_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_12_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_12_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_12_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_12_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_12_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_13_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_13_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_13_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_13_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_13_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_13_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_13_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_13_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_13_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_13_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_13_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_13_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_13_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_14_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_14_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_14_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_14_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_14_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_14_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_14_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_14_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_14_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_14_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_14_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_14_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_14_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_15_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_15_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_15_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_15_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_15_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_15_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_15_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_15_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_15_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_15_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_15_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_15_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_15_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_16_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_16_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_16_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_16_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_16_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_16_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_16_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_16_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_16_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_16_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_16_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_16_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_16_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_17_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_17_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_17_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_17_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_17_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_17_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_17_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_17_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_17_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_17_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_17_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_17_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_17_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_18_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_18_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_18_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_18_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_18_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_18_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_18_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_18_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_18_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_18_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_18_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_18_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_18_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_19_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_19_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_19_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_19_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_19_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_19_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_19_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_19_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_19_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_19_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_19_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_19_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_19_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_20_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_20_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_20_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_20_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_20_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_20_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_20_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_20_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_20_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_20_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_20_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_20_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_20_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_21_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_21_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_21_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_21_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_21_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_21_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_21_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_21_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_21_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_21_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_21_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_21_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_21_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_22_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_22_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_22_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_22_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_22_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_22_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_22_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_22_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_22_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_22_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_22_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_22_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_22_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_23_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_23_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_23_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_23_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_23_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_23_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_23_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_23_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_23_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_23_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_23_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_23_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_23_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_24_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_24_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_24_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_24_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_24_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_24_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_24_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_24_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_24_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_24_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_24_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_24_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_24_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_25_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_25_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_25_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_25_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_25_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_25_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_25_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_25_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_25_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_25_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_25_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_25_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_25_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_26_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_26_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_26_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_26_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_26_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_26_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_26_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_26_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_26_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_26_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_26_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_26_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_26_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_27_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_27_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_27_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_27_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_27_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_27_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_27_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_27_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_27_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_27_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_27_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_27_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_27_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_28_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_28_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_28_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_28_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_28_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_28_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_28_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_28_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_28_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_28_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_28_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_28_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_28_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_29_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_29_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_29_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_29_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_29_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_29_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_29_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_29_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_29_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_29_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_29_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_29_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_29_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_30_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_30_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_30_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_30_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_30_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_30_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_30_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_30_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_30_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_30_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_30_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_30_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_30_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_31_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_31_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_31_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_31_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_31_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_31_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_31_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_31_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_31_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_31_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_31_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_31_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_31_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_32_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_32_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_32_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_32_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_32_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_32_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_32_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_32_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_32_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_32_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_32_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_32_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_32_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_33_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_33_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_33_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_33_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_33_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_33_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_33_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_33_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_33_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_33_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_33_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_33_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_33_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_34_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_34_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_34_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_34_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_34_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_34_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_34_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_34_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_34_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_34_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_34_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_34_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_34_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_35_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_35_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_35_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_35_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_35_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_35_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_35_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_35_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_35_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_35_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_35_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_35_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_35_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_36_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_36_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_36_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_36_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_36_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_36_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_36_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_36_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_36_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_36_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_36_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_36_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_36_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_37_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_37_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_37_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_37_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_37_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_37_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_37_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_37_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_37_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_37_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_37_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_37_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_37_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_38_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_38_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_38_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_38_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_38_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_38_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_38_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_38_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_38_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_38_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_38_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_38_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_38_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_39_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_39_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_39_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_39_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_39_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_39_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_39_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_39_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_39_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_39_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_39_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_39_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_39_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_40_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_40_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_40_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_40_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_40_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_40_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_40_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_40_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_40_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_40_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_40_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_40_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_40_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_41_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_41_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_41_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_41_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_41_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_41_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_41_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_41_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_41_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_41_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_41_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_41_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_41_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_42_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_42_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_42_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_42_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_42_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_42_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_42_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_42_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_42_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_42_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_42_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_42_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_42_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_43_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_43_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_43_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_43_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_43_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_43_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_43_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_43_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_43_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_43_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_43_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_43_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_43_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_44_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_44_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_44_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_44_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_44_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_44_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_44_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_44_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_44_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_44_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_44_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_44_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_44_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_45_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_45_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_45_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_45_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_45_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_45_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_45_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_45_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_45_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_45_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_45_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_45_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_45_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_46_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_46_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_46_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_46_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_46_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_46_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_46_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_46_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_46_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_46_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_46_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_46_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_46_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_47_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_47_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_47_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_47_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_47_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_47_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_47_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_47_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_47_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_47_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_47_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_47_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_47_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_48_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_48_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_48_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_48_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_48_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_48_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_48_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_48_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_48_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_48_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_48_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_48_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_48_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_49_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_49_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_49_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_49_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_49_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_49_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_49_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_49_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_49_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_49_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_49_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_49_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_49_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_50_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_50_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_50_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_50_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_50_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_50_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_50_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_50_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_50_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_50_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_50_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_50_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_50_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_51_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_51_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_51_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_51_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_51_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_51_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_51_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_51_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_51_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_51_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_51_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_51_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_51_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_52_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_52_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_52_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_52_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_52_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_52_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_52_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_52_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_52_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_52_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_52_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_52_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_52_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_53_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_53_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_53_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_53_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_53_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_53_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_53_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_53_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_53_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_53_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_53_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_53_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_53_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_54_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_54_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_54_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_54_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_54_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_54_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_54_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_54_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_54_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_54_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_54_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_54_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_54_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_55_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_55_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_55_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_55_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_55_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_55_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_55_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_55_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_55_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_55_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_55_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_55_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_55_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_56_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_56_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_56_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_56_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_56_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_56_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_56_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_56_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_56_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_56_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_56_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_56_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_56_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_57_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_57_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_57_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_57_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_57_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_57_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_57_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_57_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_57_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_57_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_57_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_57_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_57_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_58_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_58_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_58_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_58_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_58_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_58_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_58_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_58_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_58_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_58_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_58_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_58_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_58_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_59_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_59_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_59_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_59_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_59_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_59_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_59_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_59_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_59_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_59_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_59_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_59_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_59_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_60_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_60_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_60_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_60_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_60_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_60_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_60_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_60_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_60_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_60_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_60_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_60_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_60_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_61_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_61_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_61_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_61_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_61_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_61_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_61_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_61_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_61_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_61_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_61_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_61_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_61_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_62_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_62_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_62_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_62_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_62_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_62_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_62_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_62_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_62_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_62_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_62_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_62_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_62_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_63_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_63_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_63_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_63_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_63_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_63_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_63_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_63_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_63_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_63_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_63_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_63_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_63_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_64_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_64_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_64_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_64_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_64_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_64_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_64_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_64_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_64_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_64_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_64_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_64_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_64_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_65_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_65_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_65_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_65_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_65_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_65_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_65_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_65_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_65_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_65_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_65_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_65_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_65_io_occupied; // @[stealNetwork.scala 23:42]
  wire  dataUnits_66_clock; // @[stealNetwork.scala 23:42]
  wire  dataUnits_66_reset; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_66_io_taskIn; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_66_io_taskOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_66_io_validIn; // @[stealNetwork.scala 23:42]
  wire  dataUnits_66_io_validOut; // @[stealNetwork.scala 23:42]
  wire  dataUnits_66_io_connSS_availableTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_66_io_connSS_availableTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_66_io_connSS_availableTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_66_io_connSS_qOutTask_ready; // @[stealNetwork.scala 23:42]
  wire  dataUnits_66_io_connSS_qOutTask_valid; // @[stealNetwork.scala 23:42]
  wire [255:0] dataUnits_66_io_connSS_qOutTask_bits; // @[stealNetwork.scala 23:42]
  wire  dataUnits_66_io_occupied; // @[stealNetwork.scala 23:42]
  wire  ctrlunits_0_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_0_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_0_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_0_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_0_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_0_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_0_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_0_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_1_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_1_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_1_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_1_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_1_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_1_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_1_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_1_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_2_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_2_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_2_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_2_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_2_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_2_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_2_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_2_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_3_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_3_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_3_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_3_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_3_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_3_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_3_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_3_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_4_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_4_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_4_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_4_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_4_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_4_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_4_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_4_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_5_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_5_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_5_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_5_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_5_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_5_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_5_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_5_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_6_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_6_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_6_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_6_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_6_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_6_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_6_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_6_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_7_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_7_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_7_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_7_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_7_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_7_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_7_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_7_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_8_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_8_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_8_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_8_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_8_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_8_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_8_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_8_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_9_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_9_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_9_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_9_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_9_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_9_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_9_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_9_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_10_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_10_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_10_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_10_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_10_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_10_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_10_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_10_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_11_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_11_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_11_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_11_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_11_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_11_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_11_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_11_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_12_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_12_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_12_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_12_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_12_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_12_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_12_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_12_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_13_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_13_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_13_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_13_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_13_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_13_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_13_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_13_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_14_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_14_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_14_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_14_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_14_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_14_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_14_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_14_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_15_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_15_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_15_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_15_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_15_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_15_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_15_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_15_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_16_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_16_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_16_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_16_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_16_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_16_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_16_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_16_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_17_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_17_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_17_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_17_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_17_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_17_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_17_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_17_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_18_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_18_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_18_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_18_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_18_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_18_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_18_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_18_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_19_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_19_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_19_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_19_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_19_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_19_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_19_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_19_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_20_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_20_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_20_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_20_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_20_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_20_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_20_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_20_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_21_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_21_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_21_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_21_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_21_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_21_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_21_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_21_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_22_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_22_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_22_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_22_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_22_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_22_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_22_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_22_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_23_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_23_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_23_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_23_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_23_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_23_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_23_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_23_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_24_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_24_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_24_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_24_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_24_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_24_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_24_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_24_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_25_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_25_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_25_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_25_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_25_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_25_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_25_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_25_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_26_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_26_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_26_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_26_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_26_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_26_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_26_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_26_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_27_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_27_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_27_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_27_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_27_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_27_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_27_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_27_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_28_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_28_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_28_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_28_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_28_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_28_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_28_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_28_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_29_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_29_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_29_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_29_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_29_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_29_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_29_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_29_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_30_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_30_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_30_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_30_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_30_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_30_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_30_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_30_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_31_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_31_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_31_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_31_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_31_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_31_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_31_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_31_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_32_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_32_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_32_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_32_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_32_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_32_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_32_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_32_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_33_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_33_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_33_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_33_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_33_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_33_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_33_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_33_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_34_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_34_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_34_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_34_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_34_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_34_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_34_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_34_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_35_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_35_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_35_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_35_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_35_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_35_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_35_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_35_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_36_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_36_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_36_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_36_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_36_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_36_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_36_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_36_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_37_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_37_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_37_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_37_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_37_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_37_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_37_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_37_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_38_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_38_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_38_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_38_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_38_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_38_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_38_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_38_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_39_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_39_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_39_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_39_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_39_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_39_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_39_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_39_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_40_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_40_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_40_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_40_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_40_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_40_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_40_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_40_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_41_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_41_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_41_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_41_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_41_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_41_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_41_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_41_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_42_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_42_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_42_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_42_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_42_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_42_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_42_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_42_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_43_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_43_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_43_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_43_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_43_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_43_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_43_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_43_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_44_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_44_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_44_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_44_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_44_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_44_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_44_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_44_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_45_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_45_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_45_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_45_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_45_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_45_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_45_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_45_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_46_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_46_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_46_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_46_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_46_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_46_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_46_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_46_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_47_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_47_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_47_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_47_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_47_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_47_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_47_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_47_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_48_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_48_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_48_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_48_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_48_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_48_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_48_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_48_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_49_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_49_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_49_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_49_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_49_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_49_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_49_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_49_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_50_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_50_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_50_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_50_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_50_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_50_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_50_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_50_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_51_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_51_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_51_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_51_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_51_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_51_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_51_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_51_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_52_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_52_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_52_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_52_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_52_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_52_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_52_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_52_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_53_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_53_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_53_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_53_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_53_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_53_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_53_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_53_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_54_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_54_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_54_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_54_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_54_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_54_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_54_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_54_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_55_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_55_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_55_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_55_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_55_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_55_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_55_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_55_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_56_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_56_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_56_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_56_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_56_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_56_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_56_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_56_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_57_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_57_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_57_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_57_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_57_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_57_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_57_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_57_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_58_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_58_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_58_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_58_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_58_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_58_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_58_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_58_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_59_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_59_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_59_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_59_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_59_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_59_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_59_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_59_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_60_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_60_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_60_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_60_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_60_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_60_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_60_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_60_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_61_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_61_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_61_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_61_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_61_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_61_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_61_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_61_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_62_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_62_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_62_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_62_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_62_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_62_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_62_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_62_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_63_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_63_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_63_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_63_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_63_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_63_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_63_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_63_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_64_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_64_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_64_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_64_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_64_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_64_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_64_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_64_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_65_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_65_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_65_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_65_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_65_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_65_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_65_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_65_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_66_clock; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_66_reset; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_66_io_reqTaskIn; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_66_io_reqTaskOut; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_66_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_66_io_connSS_serveStealReq_valid; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_66_io_connSS_stealReq_ready; // @[stealNetwork.scala 25:42]
  wire  ctrlunits_66_io_connSS_stealReq_valid; // @[stealNetwork.scala 25:42]
  stealNetworkDataUnit dataUnits_0 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_0_clock),
    .reset(dataUnits_0_reset),
    .io_taskIn(dataUnits_0_io_taskIn),
    .io_taskOut(dataUnits_0_io_taskOut),
    .io_validIn(dataUnits_0_io_validIn),
    .io_validOut(dataUnits_0_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_0_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_0_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_0_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_0_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_0_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_0_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_0_io_occupied)
  );
  stealNetworkDataUnit dataUnits_1 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_1_clock),
    .reset(dataUnits_1_reset),
    .io_taskIn(dataUnits_1_io_taskIn),
    .io_taskOut(dataUnits_1_io_taskOut),
    .io_validIn(dataUnits_1_io_validIn),
    .io_validOut(dataUnits_1_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_1_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_1_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_1_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_1_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_1_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_1_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_1_io_occupied)
  );
  stealNetworkDataUnit dataUnits_2 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_2_clock),
    .reset(dataUnits_2_reset),
    .io_taskIn(dataUnits_2_io_taskIn),
    .io_taskOut(dataUnits_2_io_taskOut),
    .io_validIn(dataUnits_2_io_validIn),
    .io_validOut(dataUnits_2_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_2_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_2_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_2_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_2_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_2_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_2_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_2_io_occupied)
  );
  stealNetworkDataUnit dataUnits_3 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_3_clock),
    .reset(dataUnits_3_reset),
    .io_taskIn(dataUnits_3_io_taskIn),
    .io_taskOut(dataUnits_3_io_taskOut),
    .io_validIn(dataUnits_3_io_validIn),
    .io_validOut(dataUnits_3_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_3_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_3_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_3_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_3_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_3_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_3_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_3_io_occupied)
  );
  stealNetworkDataUnit dataUnits_4 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_4_clock),
    .reset(dataUnits_4_reset),
    .io_taskIn(dataUnits_4_io_taskIn),
    .io_taskOut(dataUnits_4_io_taskOut),
    .io_validIn(dataUnits_4_io_validIn),
    .io_validOut(dataUnits_4_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_4_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_4_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_4_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_4_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_4_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_4_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_4_io_occupied)
  );
  stealNetworkDataUnit dataUnits_5 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_5_clock),
    .reset(dataUnits_5_reset),
    .io_taskIn(dataUnits_5_io_taskIn),
    .io_taskOut(dataUnits_5_io_taskOut),
    .io_validIn(dataUnits_5_io_validIn),
    .io_validOut(dataUnits_5_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_5_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_5_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_5_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_5_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_5_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_5_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_5_io_occupied)
  );
  stealNetworkDataUnit dataUnits_6 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_6_clock),
    .reset(dataUnits_6_reset),
    .io_taskIn(dataUnits_6_io_taskIn),
    .io_taskOut(dataUnits_6_io_taskOut),
    .io_validIn(dataUnits_6_io_validIn),
    .io_validOut(dataUnits_6_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_6_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_6_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_6_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_6_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_6_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_6_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_6_io_occupied)
  );
  stealNetworkDataUnit dataUnits_7 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_7_clock),
    .reset(dataUnits_7_reset),
    .io_taskIn(dataUnits_7_io_taskIn),
    .io_taskOut(dataUnits_7_io_taskOut),
    .io_validIn(dataUnits_7_io_validIn),
    .io_validOut(dataUnits_7_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_7_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_7_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_7_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_7_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_7_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_7_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_7_io_occupied)
  );
  stealNetworkDataUnit dataUnits_8 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_8_clock),
    .reset(dataUnits_8_reset),
    .io_taskIn(dataUnits_8_io_taskIn),
    .io_taskOut(dataUnits_8_io_taskOut),
    .io_validIn(dataUnits_8_io_validIn),
    .io_validOut(dataUnits_8_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_8_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_8_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_8_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_8_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_8_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_8_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_8_io_occupied)
  );
  stealNetworkDataUnit dataUnits_9 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_9_clock),
    .reset(dataUnits_9_reset),
    .io_taskIn(dataUnits_9_io_taskIn),
    .io_taskOut(dataUnits_9_io_taskOut),
    .io_validIn(dataUnits_9_io_validIn),
    .io_validOut(dataUnits_9_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_9_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_9_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_9_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_9_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_9_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_9_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_9_io_occupied)
  );
  stealNetworkDataUnit dataUnits_10 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_10_clock),
    .reset(dataUnits_10_reset),
    .io_taskIn(dataUnits_10_io_taskIn),
    .io_taskOut(dataUnits_10_io_taskOut),
    .io_validIn(dataUnits_10_io_validIn),
    .io_validOut(dataUnits_10_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_10_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_10_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_10_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_10_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_10_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_10_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_10_io_occupied)
  );
  stealNetworkDataUnit dataUnits_11 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_11_clock),
    .reset(dataUnits_11_reset),
    .io_taskIn(dataUnits_11_io_taskIn),
    .io_taskOut(dataUnits_11_io_taskOut),
    .io_validIn(dataUnits_11_io_validIn),
    .io_validOut(dataUnits_11_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_11_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_11_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_11_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_11_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_11_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_11_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_11_io_occupied)
  );
  stealNetworkDataUnit dataUnits_12 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_12_clock),
    .reset(dataUnits_12_reset),
    .io_taskIn(dataUnits_12_io_taskIn),
    .io_taskOut(dataUnits_12_io_taskOut),
    .io_validIn(dataUnits_12_io_validIn),
    .io_validOut(dataUnits_12_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_12_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_12_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_12_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_12_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_12_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_12_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_12_io_occupied)
  );
  stealNetworkDataUnit dataUnits_13 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_13_clock),
    .reset(dataUnits_13_reset),
    .io_taskIn(dataUnits_13_io_taskIn),
    .io_taskOut(dataUnits_13_io_taskOut),
    .io_validIn(dataUnits_13_io_validIn),
    .io_validOut(dataUnits_13_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_13_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_13_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_13_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_13_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_13_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_13_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_13_io_occupied)
  );
  stealNetworkDataUnit dataUnits_14 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_14_clock),
    .reset(dataUnits_14_reset),
    .io_taskIn(dataUnits_14_io_taskIn),
    .io_taskOut(dataUnits_14_io_taskOut),
    .io_validIn(dataUnits_14_io_validIn),
    .io_validOut(dataUnits_14_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_14_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_14_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_14_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_14_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_14_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_14_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_14_io_occupied)
  );
  stealNetworkDataUnit dataUnits_15 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_15_clock),
    .reset(dataUnits_15_reset),
    .io_taskIn(dataUnits_15_io_taskIn),
    .io_taskOut(dataUnits_15_io_taskOut),
    .io_validIn(dataUnits_15_io_validIn),
    .io_validOut(dataUnits_15_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_15_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_15_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_15_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_15_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_15_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_15_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_15_io_occupied)
  );
  stealNetworkDataUnit dataUnits_16 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_16_clock),
    .reset(dataUnits_16_reset),
    .io_taskIn(dataUnits_16_io_taskIn),
    .io_taskOut(dataUnits_16_io_taskOut),
    .io_validIn(dataUnits_16_io_validIn),
    .io_validOut(dataUnits_16_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_16_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_16_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_16_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_16_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_16_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_16_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_16_io_occupied)
  );
  stealNetworkDataUnit dataUnits_17 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_17_clock),
    .reset(dataUnits_17_reset),
    .io_taskIn(dataUnits_17_io_taskIn),
    .io_taskOut(dataUnits_17_io_taskOut),
    .io_validIn(dataUnits_17_io_validIn),
    .io_validOut(dataUnits_17_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_17_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_17_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_17_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_17_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_17_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_17_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_17_io_occupied)
  );
  stealNetworkDataUnit dataUnits_18 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_18_clock),
    .reset(dataUnits_18_reset),
    .io_taskIn(dataUnits_18_io_taskIn),
    .io_taskOut(dataUnits_18_io_taskOut),
    .io_validIn(dataUnits_18_io_validIn),
    .io_validOut(dataUnits_18_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_18_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_18_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_18_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_18_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_18_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_18_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_18_io_occupied)
  );
  stealNetworkDataUnit dataUnits_19 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_19_clock),
    .reset(dataUnits_19_reset),
    .io_taskIn(dataUnits_19_io_taskIn),
    .io_taskOut(dataUnits_19_io_taskOut),
    .io_validIn(dataUnits_19_io_validIn),
    .io_validOut(dataUnits_19_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_19_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_19_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_19_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_19_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_19_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_19_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_19_io_occupied)
  );
  stealNetworkDataUnit dataUnits_20 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_20_clock),
    .reset(dataUnits_20_reset),
    .io_taskIn(dataUnits_20_io_taskIn),
    .io_taskOut(dataUnits_20_io_taskOut),
    .io_validIn(dataUnits_20_io_validIn),
    .io_validOut(dataUnits_20_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_20_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_20_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_20_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_20_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_20_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_20_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_20_io_occupied)
  );
  stealNetworkDataUnit dataUnits_21 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_21_clock),
    .reset(dataUnits_21_reset),
    .io_taskIn(dataUnits_21_io_taskIn),
    .io_taskOut(dataUnits_21_io_taskOut),
    .io_validIn(dataUnits_21_io_validIn),
    .io_validOut(dataUnits_21_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_21_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_21_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_21_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_21_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_21_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_21_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_21_io_occupied)
  );
  stealNetworkDataUnit dataUnits_22 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_22_clock),
    .reset(dataUnits_22_reset),
    .io_taskIn(dataUnits_22_io_taskIn),
    .io_taskOut(dataUnits_22_io_taskOut),
    .io_validIn(dataUnits_22_io_validIn),
    .io_validOut(dataUnits_22_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_22_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_22_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_22_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_22_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_22_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_22_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_22_io_occupied)
  );
  stealNetworkDataUnit dataUnits_23 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_23_clock),
    .reset(dataUnits_23_reset),
    .io_taskIn(dataUnits_23_io_taskIn),
    .io_taskOut(dataUnits_23_io_taskOut),
    .io_validIn(dataUnits_23_io_validIn),
    .io_validOut(dataUnits_23_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_23_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_23_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_23_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_23_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_23_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_23_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_23_io_occupied)
  );
  stealNetworkDataUnit dataUnits_24 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_24_clock),
    .reset(dataUnits_24_reset),
    .io_taskIn(dataUnits_24_io_taskIn),
    .io_taskOut(dataUnits_24_io_taskOut),
    .io_validIn(dataUnits_24_io_validIn),
    .io_validOut(dataUnits_24_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_24_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_24_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_24_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_24_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_24_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_24_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_24_io_occupied)
  );
  stealNetworkDataUnit dataUnits_25 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_25_clock),
    .reset(dataUnits_25_reset),
    .io_taskIn(dataUnits_25_io_taskIn),
    .io_taskOut(dataUnits_25_io_taskOut),
    .io_validIn(dataUnits_25_io_validIn),
    .io_validOut(dataUnits_25_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_25_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_25_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_25_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_25_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_25_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_25_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_25_io_occupied)
  );
  stealNetworkDataUnit dataUnits_26 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_26_clock),
    .reset(dataUnits_26_reset),
    .io_taskIn(dataUnits_26_io_taskIn),
    .io_taskOut(dataUnits_26_io_taskOut),
    .io_validIn(dataUnits_26_io_validIn),
    .io_validOut(dataUnits_26_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_26_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_26_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_26_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_26_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_26_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_26_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_26_io_occupied)
  );
  stealNetworkDataUnit dataUnits_27 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_27_clock),
    .reset(dataUnits_27_reset),
    .io_taskIn(dataUnits_27_io_taskIn),
    .io_taskOut(dataUnits_27_io_taskOut),
    .io_validIn(dataUnits_27_io_validIn),
    .io_validOut(dataUnits_27_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_27_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_27_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_27_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_27_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_27_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_27_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_27_io_occupied)
  );
  stealNetworkDataUnit dataUnits_28 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_28_clock),
    .reset(dataUnits_28_reset),
    .io_taskIn(dataUnits_28_io_taskIn),
    .io_taskOut(dataUnits_28_io_taskOut),
    .io_validIn(dataUnits_28_io_validIn),
    .io_validOut(dataUnits_28_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_28_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_28_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_28_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_28_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_28_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_28_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_28_io_occupied)
  );
  stealNetworkDataUnit dataUnits_29 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_29_clock),
    .reset(dataUnits_29_reset),
    .io_taskIn(dataUnits_29_io_taskIn),
    .io_taskOut(dataUnits_29_io_taskOut),
    .io_validIn(dataUnits_29_io_validIn),
    .io_validOut(dataUnits_29_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_29_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_29_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_29_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_29_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_29_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_29_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_29_io_occupied)
  );
  stealNetworkDataUnit dataUnits_30 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_30_clock),
    .reset(dataUnits_30_reset),
    .io_taskIn(dataUnits_30_io_taskIn),
    .io_taskOut(dataUnits_30_io_taskOut),
    .io_validIn(dataUnits_30_io_validIn),
    .io_validOut(dataUnits_30_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_30_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_30_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_30_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_30_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_30_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_30_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_30_io_occupied)
  );
  stealNetworkDataUnit dataUnits_31 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_31_clock),
    .reset(dataUnits_31_reset),
    .io_taskIn(dataUnits_31_io_taskIn),
    .io_taskOut(dataUnits_31_io_taskOut),
    .io_validIn(dataUnits_31_io_validIn),
    .io_validOut(dataUnits_31_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_31_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_31_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_31_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_31_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_31_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_31_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_31_io_occupied)
  );
  stealNetworkDataUnit dataUnits_32 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_32_clock),
    .reset(dataUnits_32_reset),
    .io_taskIn(dataUnits_32_io_taskIn),
    .io_taskOut(dataUnits_32_io_taskOut),
    .io_validIn(dataUnits_32_io_validIn),
    .io_validOut(dataUnits_32_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_32_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_32_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_32_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_32_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_32_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_32_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_32_io_occupied)
  );
  stealNetworkDataUnit dataUnits_33 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_33_clock),
    .reset(dataUnits_33_reset),
    .io_taskIn(dataUnits_33_io_taskIn),
    .io_taskOut(dataUnits_33_io_taskOut),
    .io_validIn(dataUnits_33_io_validIn),
    .io_validOut(dataUnits_33_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_33_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_33_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_33_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_33_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_33_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_33_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_33_io_occupied)
  );
  stealNetworkDataUnit dataUnits_34 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_34_clock),
    .reset(dataUnits_34_reset),
    .io_taskIn(dataUnits_34_io_taskIn),
    .io_taskOut(dataUnits_34_io_taskOut),
    .io_validIn(dataUnits_34_io_validIn),
    .io_validOut(dataUnits_34_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_34_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_34_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_34_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_34_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_34_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_34_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_34_io_occupied)
  );
  stealNetworkDataUnit dataUnits_35 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_35_clock),
    .reset(dataUnits_35_reset),
    .io_taskIn(dataUnits_35_io_taskIn),
    .io_taskOut(dataUnits_35_io_taskOut),
    .io_validIn(dataUnits_35_io_validIn),
    .io_validOut(dataUnits_35_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_35_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_35_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_35_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_35_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_35_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_35_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_35_io_occupied)
  );
  stealNetworkDataUnit dataUnits_36 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_36_clock),
    .reset(dataUnits_36_reset),
    .io_taskIn(dataUnits_36_io_taskIn),
    .io_taskOut(dataUnits_36_io_taskOut),
    .io_validIn(dataUnits_36_io_validIn),
    .io_validOut(dataUnits_36_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_36_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_36_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_36_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_36_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_36_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_36_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_36_io_occupied)
  );
  stealNetworkDataUnit dataUnits_37 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_37_clock),
    .reset(dataUnits_37_reset),
    .io_taskIn(dataUnits_37_io_taskIn),
    .io_taskOut(dataUnits_37_io_taskOut),
    .io_validIn(dataUnits_37_io_validIn),
    .io_validOut(dataUnits_37_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_37_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_37_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_37_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_37_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_37_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_37_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_37_io_occupied)
  );
  stealNetworkDataUnit dataUnits_38 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_38_clock),
    .reset(dataUnits_38_reset),
    .io_taskIn(dataUnits_38_io_taskIn),
    .io_taskOut(dataUnits_38_io_taskOut),
    .io_validIn(dataUnits_38_io_validIn),
    .io_validOut(dataUnits_38_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_38_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_38_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_38_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_38_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_38_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_38_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_38_io_occupied)
  );
  stealNetworkDataUnit dataUnits_39 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_39_clock),
    .reset(dataUnits_39_reset),
    .io_taskIn(dataUnits_39_io_taskIn),
    .io_taskOut(dataUnits_39_io_taskOut),
    .io_validIn(dataUnits_39_io_validIn),
    .io_validOut(dataUnits_39_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_39_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_39_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_39_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_39_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_39_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_39_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_39_io_occupied)
  );
  stealNetworkDataUnit dataUnits_40 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_40_clock),
    .reset(dataUnits_40_reset),
    .io_taskIn(dataUnits_40_io_taskIn),
    .io_taskOut(dataUnits_40_io_taskOut),
    .io_validIn(dataUnits_40_io_validIn),
    .io_validOut(dataUnits_40_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_40_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_40_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_40_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_40_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_40_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_40_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_40_io_occupied)
  );
  stealNetworkDataUnit dataUnits_41 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_41_clock),
    .reset(dataUnits_41_reset),
    .io_taskIn(dataUnits_41_io_taskIn),
    .io_taskOut(dataUnits_41_io_taskOut),
    .io_validIn(dataUnits_41_io_validIn),
    .io_validOut(dataUnits_41_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_41_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_41_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_41_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_41_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_41_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_41_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_41_io_occupied)
  );
  stealNetworkDataUnit dataUnits_42 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_42_clock),
    .reset(dataUnits_42_reset),
    .io_taskIn(dataUnits_42_io_taskIn),
    .io_taskOut(dataUnits_42_io_taskOut),
    .io_validIn(dataUnits_42_io_validIn),
    .io_validOut(dataUnits_42_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_42_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_42_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_42_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_42_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_42_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_42_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_42_io_occupied)
  );
  stealNetworkDataUnit dataUnits_43 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_43_clock),
    .reset(dataUnits_43_reset),
    .io_taskIn(dataUnits_43_io_taskIn),
    .io_taskOut(dataUnits_43_io_taskOut),
    .io_validIn(dataUnits_43_io_validIn),
    .io_validOut(dataUnits_43_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_43_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_43_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_43_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_43_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_43_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_43_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_43_io_occupied)
  );
  stealNetworkDataUnit dataUnits_44 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_44_clock),
    .reset(dataUnits_44_reset),
    .io_taskIn(dataUnits_44_io_taskIn),
    .io_taskOut(dataUnits_44_io_taskOut),
    .io_validIn(dataUnits_44_io_validIn),
    .io_validOut(dataUnits_44_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_44_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_44_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_44_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_44_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_44_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_44_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_44_io_occupied)
  );
  stealNetworkDataUnit dataUnits_45 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_45_clock),
    .reset(dataUnits_45_reset),
    .io_taskIn(dataUnits_45_io_taskIn),
    .io_taskOut(dataUnits_45_io_taskOut),
    .io_validIn(dataUnits_45_io_validIn),
    .io_validOut(dataUnits_45_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_45_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_45_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_45_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_45_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_45_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_45_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_45_io_occupied)
  );
  stealNetworkDataUnit dataUnits_46 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_46_clock),
    .reset(dataUnits_46_reset),
    .io_taskIn(dataUnits_46_io_taskIn),
    .io_taskOut(dataUnits_46_io_taskOut),
    .io_validIn(dataUnits_46_io_validIn),
    .io_validOut(dataUnits_46_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_46_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_46_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_46_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_46_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_46_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_46_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_46_io_occupied)
  );
  stealNetworkDataUnit dataUnits_47 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_47_clock),
    .reset(dataUnits_47_reset),
    .io_taskIn(dataUnits_47_io_taskIn),
    .io_taskOut(dataUnits_47_io_taskOut),
    .io_validIn(dataUnits_47_io_validIn),
    .io_validOut(dataUnits_47_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_47_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_47_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_47_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_47_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_47_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_47_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_47_io_occupied)
  );
  stealNetworkDataUnit dataUnits_48 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_48_clock),
    .reset(dataUnits_48_reset),
    .io_taskIn(dataUnits_48_io_taskIn),
    .io_taskOut(dataUnits_48_io_taskOut),
    .io_validIn(dataUnits_48_io_validIn),
    .io_validOut(dataUnits_48_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_48_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_48_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_48_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_48_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_48_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_48_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_48_io_occupied)
  );
  stealNetworkDataUnit dataUnits_49 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_49_clock),
    .reset(dataUnits_49_reset),
    .io_taskIn(dataUnits_49_io_taskIn),
    .io_taskOut(dataUnits_49_io_taskOut),
    .io_validIn(dataUnits_49_io_validIn),
    .io_validOut(dataUnits_49_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_49_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_49_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_49_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_49_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_49_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_49_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_49_io_occupied)
  );
  stealNetworkDataUnit dataUnits_50 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_50_clock),
    .reset(dataUnits_50_reset),
    .io_taskIn(dataUnits_50_io_taskIn),
    .io_taskOut(dataUnits_50_io_taskOut),
    .io_validIn(dataUnits_50_io_validIn),
    .io_validOut(dataUnits_50_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_50_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_50_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_50_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_50_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_50_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_50_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_50_io_occupied)
  );
  stealNetworkDataUnit dataUnits_51 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_51_clock),
    .reset(dataUnits_51_reset),
    .io_taskIn(dataUnits_51_io_taskIn),
    .io_taskOut(dataUnits_51_io_taskOut),
    .io_validIn(dataUnits_51_io_validIn),
    .io_validOut(dataUnits_51_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_51_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_51_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_51_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_51_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_51_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_51_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_51_io_occupied)
  );
  stealNetworkDataUnit dataUnits_52 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_52_clock),
    .reset(dataUnits_52_reset),
    .io_taskIn(dataUnits_52_io_taskIn),
    .io_taskOut(dataUnits_52_io_taskOut),
    .io_validIn(dataUnits_52_io_validIn),
    .io_validOut(dataUnits_52_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_52_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_52_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_52_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_52_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_52_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_52_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_52_io_occupied)
  );
  stealNetworkDataUnit dataUnits_53 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_53_clock),
    .reset(dataUnits_53_reset),
    .io_taskIn(dataUnits_53_io_taskIn),
    .io_taskOut(dataUnits_53_io_taskOut),
    .io_validIn(dataUnits_53_io_validIn),
    .io_validOut(dataUnits_53_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_53_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_53_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_53_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_53_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_53_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_53_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_53_io_occupied)
  );
  stealNetworkDataUnit dataUnits_54 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_54_clock),
    .reset(dataUnits_54_reset),
    .io_taskIn(dataUnits_54_io_taskIn),
    .io_taskOut(dataUnits_54_io_taskOut),
    .io_validIn(dataUnits_54_io_validIn),
    .io_validOut(dataUnits_54_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_54_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_54_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_54_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_54_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_54_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_54_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_54_io_occupied)
  );
  stealNetworkDataUnit dataUnits_55 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_55_clock),
    .reset(dataUnits_55_reset),
    .io_taskIn(dataUnits_55_io_taskIn),
    .io_taskOut(dataUnits_55_io_taskOut),
    .io_validIn(dataUnits_55_io_validIn),
    .io_validOut(dataUnits_55_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_55_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_55_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_55_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_55_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_55_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_55_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_55_io_occupied)
  );
  stealNetworkDataUnit dataUnits_56 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_56_clock),
    .reset(dataUnits_56_reset),
    .io_taskIn(dataUnits_56_io_taskIn),
    .io_taskOut(dataUnits_56_io_taskOut),
    .io_validIn(dataUnits_56_io_validIn),
    .io_validOut(dataUnits_56_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_56_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_56_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_56_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_56_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_56_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_56_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_56_io_occupied)
  );
  stealNetworkDataUnit dataUnits_57 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_57_clock),
    .reset(dataUnits_57_reset),
    .io_taskIn(dataUnits_57_io_taskIn),
    .io_taskOut(dataUnits_57_io_taskOut),
    .io_validIn(dataUnits_57_io_validIn),
    .io_validOut(dataUnits_57_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_57_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_57_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_57_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_57_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_57_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_57_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_57_io_occupied)
  );
  stealNetworkDataUnit dataUnits_58 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_58_clock),
    .reset(dataUnits_58_reset),
    .io_taskIn(dataUnits_58_io_taskIn),
    .io_taskOut(dataUnits_58_io_taskOut),
    .io_validIn(dataUnits_58_io_validIn),
    .io_validOut(dataUnits_58_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_58_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_58_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_58_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_58_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_58_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_58_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_58_io_occupied)
  );
  stealNetworkDataUnit dataUnits_59 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_59_clock),
    .reset(dataUnits_59_reset),
    .io_taskIn(dataUnits_59_io_taskIn),
    .io_taskOut(dataUnits_59_io_taskOut),
    .io_validIn(dataUnits_59_io_validIn),
    .io_validOut(dataUnits_59_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_59_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_59_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_59_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_59_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_59_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_59_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_59_io_occupied)
  );
  stealNetworkDataUnit dataUnits_60 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_60_clock),
    .reset(dataUnits_60_reset),
    .io_taskIn(dataUnits_60_io_taskIn),
    .io_taskOut(dataUnits_60_io_taskOut),
    .io_validIn(dataUnits_60_io_validIn),
    .io_validOut(dataUnits_60_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_60_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_60_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_60_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_60_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_60_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_60_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_60_io_occupied)
  );
  stealNetworkDataUnit dataUnits_61 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_61_clock),
    .reset(dataUnits_61_reset),
    .io_taskIn(dataUnits_61_io_taskIn),
    .io_taskOut(dataUnits_61_io_taskOut),
    .io_validIn(dataUnits_61_io_validIn),
    .io_validOut(dataUnits_61_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_61_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_61_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_61_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_61_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_61_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_61_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_61_io_occupied)
  );
  stealNetworkDataUnit dataUnits_62 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_62_clock),
    .reset(dataUnits_62_reset),
    .io_taskIn(dataUnits_62_io_taskIn),
    .io_taskOut(dataUnits_62_io_taskOut),
    .io_validIn(dataUnits_62_io_validIn),
    .io_validOut(dataUnits_62_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_62_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_62_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_62_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_62_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_62_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_62_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_62_io_occupied)
  );
  stealNetworkDataUnit dataUnits_63 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_63_clock),
    .reset(dataUnits_63_reset),
    .io_taskIn(dataUnits_63_io_taskIn),
    .io_taskOut(dataUnits_63_io_taskOut),
    .io_validIn(dataUnits_63_io_validIn),
    .io_validOut(dataUnits_63_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_63_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_63_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_63_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_63_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_63_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_63_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_63_io_occupied)
  );
  stealNetworkDataUnit dataUnits_64 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_64_clock),
    .reset(dataUnits_64_reset),
    .io_taskIn(dataUnits_64_io_taskIn),
    .io_taskOut(dataUnits_64_io_taskOut),
    .io_validIn(dataUnits_64_io_validIn),
    .io_validOut(dataUnits_64_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_64_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_64_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_64_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_64_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_64_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_64_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_64_io_occupied)
  );
  stealNetworkDataUnit dataUnits_65 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_65_clock),
    .reset(dataUnits_65_reset),
    .io_taskIn(dataUnits_65_io_taskIn),
    .io_taskOut(dataUnits_65_io_taskOut),
    .io_validIn(dataUnits_65_io_validIn),
    .io_validOut(dataUnits_65_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_65_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_65_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_65_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_65_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_65_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_65_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_65_io_occupied)
  );
  stealNetworkDataUnit dataUnits_66 ( // @[stealNetwork.scala 23:42]
    .clock(dataUnits_66_clock),
    .reset(dataUnits_66_reset),
    .io_taskIn(dataUnits_66_io_taskIn),
    .io_taskOut(dataUnits_66_io_taskOut),
    .io_validIn(dataUnits_66_io_validIn),
    .io_validOut(dataUnits_66_io_validOut),
    .io_connSS_availableTask_ready(dataUnits_66_io_connSS_availableTask_ready),
    .io_connSS_availableTask_valid(dataUnits_66_io_connSS_availableTask_valid),
    .io_connSS_availableTask_bits(dataUnits_66_io_connSS_availableTask_bits),
    .io_connSS_qOutTask_ready(dataUnits_66_io_connSS_qOutTask_ready),
    .io_connSS_qOutTask_valid(dataUnits_66_io_connSS_qOutTask_valid),
    .io_connSS_qOutTask_bits(dataUnits_66_io_connSS_qOutTask_bits),
    .io_occupied(dataUnits_66_io_occupied)
  );
  stealNetworkCtrlUnit ctrlunits_0 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_0_clock),
    .reset(ctrlunits_0_reset),
    .io_reqTaskIn(ctrlunits_0_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_0_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_0_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_0_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_0_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_0_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_1 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_1_clock),
    .reset(ctrlunits_1_reset),
    .io_reqTaskIn(ctrlunits_1_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_1_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_1_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_1_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_1_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_1_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_2 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_2_clock),
    .reset(ctrlunits_2_reset),
    .io_reqTaskIn(ctrlunits_2_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_2_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_2_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_2_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_2_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_2_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_3 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_3_clock),
    .reset(ctrlunits_3_reset),
    .io_reqTaskIn(ctrlunits_3_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_3_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_3_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_3_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_3_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_3_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_4 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_4_clock),
    .reset(ctrlunits_4_reset),
    .io_reqTaskIn(ctrlunits_4_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_4_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_4_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_4_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_4_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_4_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_5 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_5_clock),
    .reset(ctrlunits_5_reset),
    .io_reqTaskIn(ctrlunits_5_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_5_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_5_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_5_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_5_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_5_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_6 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_6_clock),
    .reset(ctrlunits_6_reset),
    .io_reqTaskIn(ctrlunits_6_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_6_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_6_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_6_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_6_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_6_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_7 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_7_clock),
    .reset(ctrlunits_7_reset),
    .io_reqTaskIn(ctrlunits_7_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_7_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_7_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_7_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_7_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_7_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_8 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_8_clock),
    .reset(ctrlunits_8_reset),
    .io_reqTaskIn(ctrlunits_8_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_8_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_8_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_8_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_8_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_8_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_9 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_9_clock),
    .reset(ctrlunits_9_reset),
    .io_reqTaskIn(ctrlunits_9_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_9_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_9_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_9_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_9_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_9_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_10 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_10_clock),
    .reset(ctrlunits_10_reset),
    .io_reqTaskIn(ctrlunits_10_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_10_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_10_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_10_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_10_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_10_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_11 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_11_clock),
    .reset(ctrlunits_11_reset),
    .io_reqTaskIn(ctrlunits_11_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_11_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_11_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_11_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_11_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_11_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_12 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_12_clock),
    .reset(ctrlunits_12_reset),
    .io_reqTaskIn(ctrlunits_12_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_12_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_12_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_12_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_12_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_12_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_13 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_13_clock),
    .reset(ctrlunits_13_reset),
    .io_reqTaskIn(ctrlunits_13_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_13_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_13_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_13_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_13_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_13_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_14 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_14_clock),
    .reset(ctrlunits_14_reset),
    .io_reqTaskIn(ctrlunits_14_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_14_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_14_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_14_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_14_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_14_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_15 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_15_clock),
    .reset(ctrlunits_15_reset),
    .io_reqTaskIn(ctrlunits_15_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_15_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_15_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_15_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_15_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_15_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_16 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_16_clock),
    .reset(ctrlunits_16_reset),
    .io_reqTaskIn(ctrlunits_16_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_16_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_16_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_16_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_16_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_16_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_17 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_17_clock),
    .reset(ctrlunits_17_reset),
    .io_reqTaskIn(ctrlunits_17_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_17_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_17_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_17_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_17_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_17_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_18 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_18_clock),
    .reset(ctrlunits_18_reset),
    .io_reqTaskIn(ctrlunits_18_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_18_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_18_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_18_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_18_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_18_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_19 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_19_clock),
    .reset(ctrlunits_19_reset),
    .io_reqTaskIn(ctrlunits_19_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_19_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_19_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_19_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_19_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_19_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_20 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_20_clock),
    .reset(ctrlunits_20_reset),
    .io_reqTaskIn(ctrlunits_20_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_20_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_20_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_20_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_20_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_20_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_21 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_21_clock),
    .reset(ctrlunits_21_reset),
    .io_reqTaskIn(ctrlunits_21_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_21_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_21_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_21_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_21_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_21_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_22 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_22_clock),
    .reset(ctrlunits_22_reset),
    .io_reqTaskIn(ctrlunits_22_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_22_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_22_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_22_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_22_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_22_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_23 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_23_clock),
    .reset(ctrlunits_23_reset),
    .io_reqTaskIn(ctrlunits_23_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_23_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_23_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_23_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_23_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_23_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_24 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_24_clock),
    .reset(ctrlunits_24_reset),
    .io_reqTaskIn(ctrlunits_24_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_24_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_24_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_24_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_24_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_24_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_25 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_25_clock),
    .reset(ctrlunits_25_reset),
    .io_reqTaskIn(ctrlunits_25_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_25_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_25_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_25_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_25_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_25_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_26 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_26_clock),
    .reset(ctrlunits_26_reset),
    .io_reqTaskIn(ctrlunits_26_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_26_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_26_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_26_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_26_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_26_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_27 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_27_clock),
    .reset(ctrlunits_27_reset),
    .io_reqTaskIn(ctrlunits_27_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_27_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_27_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_27_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_27_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_27_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_28 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_28_clock),
    .reset(ctrlunits_28_reset),
    .io_reqTaskIn(ctrlunits_28_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_28_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_28_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_28_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_28_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_28_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_29 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_29_clock),
    .reset(ctrlunits_29_reset),
    .io_reqTaskIn(ctrlunits_29_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_29_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_29_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_29_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_29_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_29_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_30 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_30_clock),
    .reset(ctrlunits_30_reset),
    .io_reqTaskIn(ctrlunits_30_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_30_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_30_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_30_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_30_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_30_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_31 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_31_clock),
    .reset(ctrlunits_31_reset),
    .io_reqTaskIn(ctrlunits_31_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_31_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_31_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_31_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_31_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_31_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_32 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_32_clock),
    .reset(ctrlunits_32_reset),
    .io_reqTaskIn(ctrlunits_32_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_32_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_32_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_32_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_32_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_32_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_33 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_33_clock),
    .reset(ctrlunits_33_reset),
    .io_reqTaskIn(ctrlunits_33_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_33_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_33_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_33_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_33_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_33_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_34 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_34_clock),
    .reset(ctrlunits_34_reset),
    .io_reqTaskIn(ctrlunits_34_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_34_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_34_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_34_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_34_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_34_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_35 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_35_clock),
    .reset(ctrlunits_35_reset),
    .io_reqTaskIn(ctrlunits_35_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_35_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_35_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_35_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_35_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_35_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_36 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_36_clock),
    .reset(ctrlunits_36_reset),
    .io_reqTaskIn(ctrlunits_36_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_36_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_36_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_36_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_36_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_36_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_37 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_37_clock),
    .reset(ctrlunits_37_reset),
    .io_reqTaskIn(ctrlunits_37_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_37_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_37_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_37_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_37_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_37_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_38 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_38_clock),
    .reset(ctrlunits_38_reset),
    .io_reqTaskIn(ctrlunits_38_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_38_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_38_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_38_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_38_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_38_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_39 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_39_clock),
    .reset(ctrlunits_39_reset),
    .io_reqTaskIn(ctrlunits_39_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_39_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_39_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_39_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_39_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_39_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_40 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_40_clock),
    .reset(ctrlunits_40_reset),
    .io_reqTaskIn(ctrlunits_40_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_40_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_40_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_40_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_40_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_40_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_41 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_41_clock),
    .reset(ctrlunits_41_reset),
    .io_reqTaskIn(ctrlunits_41_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_41_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_41_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_41_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_41_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_41_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_42 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_42_clock),
    .reset(ctrlunits_42_reset),
    .io_reqTaskIn(ctrlunits_42_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_42_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_42_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_42_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_42_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_42_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_43 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_43_clock),
    .reset(ctrlunits_43_reset),
    .io_reqTaskIn(ctrlunits_43_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_43_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_43_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_43_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_43_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_43_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_44 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_44_clock),
    .reset(ctrlunits_44_reset),
    .io_reqTaskIn(ctrlunits_44_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_44_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_44_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_44_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_44_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_44_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_45 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_45_clock),
    .reset(ctrlunits_45_reset),
    .io_reqTaskIn(ctrlunits_45_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_45_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_45_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_45_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_45_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_45_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_46 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_46_clock),
    .reset(ctrlunits_46_reset),
    .io_reqTaskIn(ctrlunits_46_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_46_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_46_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_46_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_46_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_46_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_47 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_47_clock),
    .reset(ctrlunits_47_reset),
    .io_reqTaskIn(ctrlunits_47_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_47_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_47_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_47_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_47_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_47_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_48 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_48_clock),
    .reset(ctrlunits_48_reset),
    .io_reqTaskIn(ctrlunits_48_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_48_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_48_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_48_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_48_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_48_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_49 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_49_clock),
    .reset(ctrlunits_49_reset),
    .io_reqTaskIn(ctrlunits_49_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_49_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_49_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_49_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_49_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_49_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_50 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_50_clock),
    .reset(ctrlunits_50_reset),
    .io_reqTaskIn(ctrlunits_50_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_50_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_50_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_50_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_50_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_50_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_51 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_51_clock),
    .reset(ctrlunits_51_reset),
    .io_reqTaskIn(ctrlunits_51_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_51_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_51_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_51_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_51_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_51_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_52 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_52_clock),
    .reset(ctrlunits_52_reset),
    .io_reqTaskIn(ctrlunits_52_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_52_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_52_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_52_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_52_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_52_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_53 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_53_clock),
    .reset(ctrlunits_53_reset),
    .io_reqTaskIn(ctrlunits_53_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_53_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_53_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_53_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_53_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_53_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_54 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_54_clock),
    .reset(ctrlunits_54_reset),
    .io_reqTaskIn(ctrlunits_54_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_54_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_54_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_54_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_54_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_54_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_55 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_55_clock),
    .reset(ctrlunits_55_reset),
    .io_reqTaskIn(ctrlunits_55_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_55_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_55_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_55_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_55_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_55_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_56 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_56_clock),
    .reset(ctrlunits_56_reset),
    .io_reqTaskIn(ctrlunits_56_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_56_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_56_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_56_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_56_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_56_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_57 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_57_clock),
    .reset(ctrlunits_57_reset),
    .io_reqTaskIn(ctrlunits_57_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_57_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_57_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_57_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_57_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_57_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_58 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_58_clock),
    .reset(ctrlunits_58_reset),
    .io_reqTaskIn(ctrlunits_58_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_58_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_58_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_58_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_58_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_58_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_59 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_59_clock),
    .reset(ctrlunits_59_reset),
    .io_reqTaskIn(ctrlunits_59_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_59_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_59_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_59_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_59_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_59_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_60 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_60_clock),
    .reset(ctrlunits_60_reset),
    .io_reqTaskIn(ctrlunits_60_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_60_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_60_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_60_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_60_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_60_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_61 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_61_clock),
    .reset(ctrlunits_61_reset),
    .io_reqTaskIn(ctrlunits_61_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_61_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_61_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_61_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_61_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_61_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_62 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_62_clock),
    .reset(ctrlunits_62_reset),
    .io_reqTaskIn(ctrlunits_62_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_62_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_62_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_62_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_62_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_62_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_63 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_63_clock),
    .reset(ctrlunits_63_reset),
    .io_reqTaskIn(ctrlunits_63_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_63_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_63_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_63_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_63_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_63_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_64 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_64_clock),
    .reset(ctrlunits_64_reset),
    .io_reqTaskIn(ctrlunits_64_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_64_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_64_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_64_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_64_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_64_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_65 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_65_clock),
    .reset(ctrlunits_65_reset),
    .io_reqTaskIn(ctrlunits_65_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_65_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_65_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_65_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_65_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_65_io_connSS_stealReq_valid)
  );
  stealNetworkCtrlUnit ctrlunits_66 ( // @[stealNetwork.scala 25:42]
    .clock(ctrlunits_66_clock),
    .reset(ctrlunits_66_reset),
    .io_reqTaskIn(ctrlunits_66_io_reqTaskIn),
    .io_reqTaskOut(ctrlunits_66_io_reqTaskOut),
    .io_connSS_serveStealReq_ready(ctrlunits_66_io_connSS_serveStealReq_ready),
    .io_connSS_serveStealReq_valid(ctrlunits_66_io_connSS_serveStealReq_valid),
    .io_connSS_stealReq_ready(ctrlunits_66_io_connSS_stealReq_ready),
    .io_connSS_stealReq_valid(ctrlunits_66_io_connSS_stealReq_valid)
  );
  assign io_connSS_0_ctrl_serveStealReq_ready = ctrlunits_0_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_0_data_availableTask_valid = dataUnits_0_io_connSS_availableTask_valid; // @[stealNetwork.scala 36:27]
  assign io_connSS_0_data_availableTask_bits = dataUnits_0_io_connSS_availableTask_bits; // @[stealNetwork.scala 36:27]
  assign io_connSS_0_data_qOutTask_ready = dataUnits_0_io_connSS_qOutTask_ready; // @[stealNetwork.scala 36:27]
  assign io_connSS_1_ctrl_serveStealReq_ready = ctrlunits_1_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_1_data_qOutTask_ready = dataUnits_1_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_2_ctrl_serveStealReq_ready = ctrlunits_2_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_2_data_qOutTask_ready = dataUnits_2_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_3_ctrl_serveStealReq_ready = ctrlunits_3_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_3_ctrl_stealReq_ready = ctrlunits_3_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_3_data_availableTask_valid = dataUnits_3_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_3_data_availableTask_bits = dataUnits_3_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_3_data_qOutTask_ready = dataUnits_3_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_4_ctrl_serveStealReq_ready = ctrlunits_4_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_4_ctrl_stealReq_ready = ctrlunits_4_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_4_data_availableTask_valid = dataUnits_4_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_4_data_availableTask_bits = dataUnits_4_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_4_data_qOutTask_ready = dataUnits_4_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_5_ctrl_serveStealReq_ready = ctrlunits_5_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_5_ctrl_stealReq_ready = ctrlunits_5_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_5_data_availableTask_valid = dataUnits_5_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_5_data_availableTask_bits = dataUnits_5_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_5_data_qOutTask_ready = dataUnits_5_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_6_ctrl_serveStealReq_ready = ctrlunits_6_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_6_ctrl_stealReq_ready = ctrlunits_6_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_6_data_availableTask_valid = dataUnits_6_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_6_data_availableTask_bits = dataUnits_6_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_6_data_qOutTask_ready = dataUnits_6_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_7_ctrl_serveStealReq_ready = ctrlunits_7_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_7_ctrl_stealReq_ready = ctrlunits_7_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_7_data_availableTask_valid = dataUnits_7_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_7_data_availableTask_bits = dataUnits_7_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_7_data_qOutTask_ready = dataUnits_7_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_8_ctrl_serveStealReq_ready = ctrlunits_8_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_8_ctrl_stealReq_ready = ctrlunits_8_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_8_data_availableTask_valid = dataUnits_8_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_8_data_availableTask_bits = dataUnits_8_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_8_data_qOutTask_ready = dataUnits_8_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_9_ctrl_serveStealReq_ready = ctrlunits_9_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_9_ctrl_stealReq_ready = ctrlunits_9_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_9_data_availableTask_valid = dataUnits_9_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_9_data_availableTask_bits = dataUnits_9_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_9_data_qOutTask_ready = dataUnits_9_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_10_ctrl_serveStealReq_ready = ctrlunits_10_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_10_ctrl_stealReq_ready = ctrlunits_10_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_10_data_availableTask_valid = dataUnits_10_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_10_data_availableTask_bits = dataUnits_10_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_10_data_qOutTask_ready = dataUnits_10_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_11_ctrl_serveStealReq_ready = ctrlunits_11_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_11_ctrl_stealReq_ready = ctrlunits_11_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_11_data_availableTask_valid = dataUnits_11_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_11_data_availableTask_bits = dataUnits_11_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_11_data_qOutTask_ready = dataUnits_11_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_12_ctrl_serveStealReq_ready = ctrlunits_12_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_12_ctrl_stealReq_ready = ctrlunits_12_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_12_data_availableTask_valid = dataUnits_12_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_12_data_availableTask_bits = dataUnits_12_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_12_data_qOutTask_ready = dataUnits_12_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_13_ctrl_serveStealReq_ready = ctrlunits_13_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_13_ctrl_stealReq_ready = ctrlunits_13_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_13_data_availableTask_valid = dataUnits_13_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_13_data_availableTask_bits = dataUnits_13_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_13_data_qOutTask_ready = dataUnits_13_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_14_ctrl_serveStealReq_ready = ctrlunits_14_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_14_ctrl_stealReq_ready = ctrlunits_14_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_14_data_availableTask_valid = dataUnits_14_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_14_data_availableTask_bits = dataUnits_14_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_14_data_qOutTask_ready = dataUnits_14_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_15_ctrl_serveStealReq_ready = ctrlunits_15_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_15_ctrl_stealReq_ready = ctrlunits_15_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_15_data_availableTask_valid = dataUnits_15_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_15_data_availableTask_bits = dataUnits_15_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_15_data_qOutTask_ready = dataUnits_15_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_16_ctrl_serveStealReq_ready = ctrlunits_16_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_16_ctrl_stealReq_ready = ctrlunits_16_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_16_data_availableTask_valid = dataUnits_16_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_16_data_availableTask_bits = dataUnits_16_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_16_data_qOutTask_ready = dataUnits_16_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_17_ctrl_serveStealReq_ready = ctrlunits_17_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_17_ctrl_stealReq_ready = ctrlunits_17_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_17_data_availableTask_valid = dataUnits_17_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_17_data_availableTask_bits = dataUnits_17_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_17_data_qOutTask_ready = dataUnits_17_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_18_ctrl_serveStealReq_ready = ctrlunits_18_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_18_ctrl_stealReq_ready = ctrlunits_18_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_18_data_availableTask_valid = dataUnits_18_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_18_data_availableTask_bits = dataUnits_18_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_18_data_qOutTask_ready = dataUnits_18_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_19_ctrl_serveStealReq_ready = ctrlunits_19_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_19_ctrl_stealReq_ready = ctrlunits_19_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_19_data_availableTask_valid = dataUnits_19_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_19_data_availableTask_bits = dataUnits_19_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_19_data_qOutTask_ready = dataUnits_19_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_20_ctrl_serveStealReq_ready = ctrlunits_20_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_20_ctrl_stealReq_ready = ctrlunits_20_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_20_data_availableTask_valid = dataUnits_20_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_20_data_availableTask_bits = dataUnits_20_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_20_data_qOutTask_ready = dataUnits_20_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_21_ctrl_serveStealReq_ready = ctrlunits_21_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_21_ctrl_stealReq_ready = ctrlunits_21_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_21_data_availableTask_valid = dataUnits_21_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_21_data_availableTask_bits = dataUnits_21_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_21_data_qOutTask_ready = dataUnits_21_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_22_ctrl_serveStealReq_ready = ctrlunits_22_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_22_ctrl_stealReq_ready = ctrlunits_22_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_22_data_availableTask_valid = dataUnits_22_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_22_data_availableTask_bits = dataUnits_22_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_22_data_qOutTask_ready = dataUnits_22_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_23_ctrl_serveStealReq_ready = ctrlunits_23_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_23_ctrl_stealReq_ready = ctrlunits_23_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_23_data_availableTask_valid = dataUnits_23_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_23_data_availableTask_bits = dataUnits_23_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_23_data_qOutTask_ready = dataUnits_23_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_24_ctrl_serveStealReq_ready = ctrlunits_24_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_24_ctrl_stealReq_ready = ctrlunits_24_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_24_data_availableTask_valid = dataUnits_24_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_24_data_availableTask_bits = dataUnits_24_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_24_data_qOutTask_ready = dataUnits_24_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_25_ctrl_serveStealReq_ready = ctrlunits_25_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_25_ctrl_stealReq_ready = ctrlunits_25_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_25_data_availableTask_valid = dataUnits_25_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_25_data_availableTask_bits = dataUnits_25_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_25_data_qOutTask_ready = dataUnits_25_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_26_ctrl_serveStealReq_ready = ctrlunits_26_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_26_ctrl_stealReq_ready = ctrlunits_26_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_26_data_availableTask_valid = dataUnits_26_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_26_data_availableTask_bits = dataUnits_26_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_26_data_qOutTask_ready = dataUnits_26_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_27_ctrl_serveStealReq_ready = ctrlunits_27_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_27_ctrl_stealReq_ready = ctrlunits_27_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_27_data_availableTask_valid = dataUnits_27_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_27_data_availableTask_bits = dataUnits_27_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_27_data_qOutTask_ready = dataUnits_27_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_28_ctrl_serveStealReq_ready = ctrlunits_28_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_28_ctrl_stealReq_ready = ctrlunits_28_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_28_data_availableTask_valid = dataUnits_28_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_28_data_availableTask_bits = dataUnits_28_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_28_data_qOutTask_ready = dataUnits_28_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_29_ctrl_serveStealReq_ready = ctrlunits_29_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_29_ctrl_stealReq_ready = ctrlunits_29_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_29_data_availableTask_valid = dataUnits_29_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_29_data_availableTask_bits = dataUnits_29_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_29_data_qOutTask_ready = dataUnits_29_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_30_ctrl_serveStealReq_ready = ctrlunits_30_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_30_ctrl_stealReq_ready = ctrlunits_30_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_30_data_availableTask_valid = dataUnits_30_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_30_data_availableTask_bits = dataUnits_30_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_30_data_qOutTask_ready = dataUnits_30_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_31_ctrl_serveStealReq_ready = ctrlunits_31_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_31_ctrl_stealReq_ready = ctrlunits_31_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_31_data_availableTask_valid = dataUnits_31_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_31_data_availableTask_bits = dataUnits_31_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_31_data_qOutTask_ready = dataUnits_31_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_32_ctrl_serveStealReq_ready = ctrlunits_32_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_32_ctrl_stealReq_ready = ctrlunits_32_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_32_data_availableTask_valid = dataUnits_32_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_32_data_availableTask_bits = dataUnits_32_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_32_data_qOutTask_ready = dataUnits_32_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_33_ctrl_serveStealReq_ready = ctrlunits_33_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_33_ctrl_stealReq_ready = ctrlunits_33_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_33_data_availableTask_valid = dataUnits_33_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_33_data_availableTask_bits = dataUnits_33_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_33_data_qOutTask_ready = dataUnits_33_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_34_ctrl_serveStealReq_ready = ctrlunits_34_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_34_ctrl_stealReq_ready = ctrlunits_34_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_34_data_availableTask_valid = dataUnits_34_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_34_data_availableTask_bits = dataUnits_34_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_34_data_qOutTask_ready = dataUnits_34_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_35_ctrl_serveStealReq_ready = ctrlunits_35_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_35_ctrl_stealReq_ready = ctrlunits_35_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_35_data_availableTask_valid = dataUnits_35_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_35_data_availableTask_bits = dataUnits_35_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_35_data_qOutTask_ready = dataUnits_35_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_36_ctrl_serveStealReq_ready = ctrlunits_36_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_36_ctrl_stealReq_ready = ctrlunits_36_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_36_data_availableTask_valid = dataUnits_36_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_36_data_availableTask_bits = dataUnits_36_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_36_data_qOutTask_ready = dataUnits_36_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_37_ctrl_serveStealReq_ready = ctrlunits_37_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_37_ctrl_stealReq_ready = ctrlunits_37_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_37_data_availableTask_valid = dataUnits_37_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_37_data_availableTask_bits = dataUnits_37_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_37_data_qOutTask_ready = dataUnits_37_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_38_ctrl_serveStealReq_ready = ctrlunits_38_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_38_ctrl_stealReq_ready = ctrlunits_38_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_38_data_availableTask_valid = dataUnits_38_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_38_data_availableTask_bits = dataUnits_38_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_38_data_qOutTask_ready = dataUnits_38_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_39_ctrl_serveStealReq_ready = ctrlunits_39_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_39_ctrl_stealReq_ready = ctrlunits_39_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_39_data_availableTask_valid = dataUnits_39_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_39_data_availableTask_bits = dataUnits_39_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_39_data_qOutTask_ready = dataUnits_39_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_40_ctrl_serveStealReq_ready = ctrlunits_40_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_40_ctrl_stealReq_ready = ctrlunits_40_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_40_data_availableTask_valid = dataUnits_40_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_40_data_availableTask_bits = dataUnits_40_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_40_data_qOutTask_ready = dataUnits_40_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_41_ctrl_serveStealReq_ready = ctrlunits_41_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_41_ctrl_stealReq_ready = ctrlunits_41_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_41_data_availableTask_valid = dataUnits_41_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_41_data_availableTask_bits = dataUnits_41_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_41_data_qOutTask_ready = dataUnits_41_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_42_ctrl_serveStealReq_ready = ctrlunits_42_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_42_ctrl_stealReq_ready = ctrlunits_42_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_42_data_availableTask_valid = dataUnits_42_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_42_data_availableTask_bits = dataUnits_42_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_42_data_qOutTask_ready = dataUnits_42_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_43_ctrl_serveStealReq_ready = ctrlunits_43_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_43_ctrl_stealReq_ready = ctrlunits_43_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_43_data_availableTask_valid = dataUnits_43_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_43_data_availableTask_bits = dataUnits_43_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_43_data_qOutTask_ready = dataUnits_43_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_44_ctrl_serveStealReq_ready = ctrlunits_44_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_44_ctrl_stealReq_ready = ctrlunits_44_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_44_data_availableTask_valid = dataUnits_44_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_44_data_availableTask_bits = dataUnits_44_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_44_data_qOutTask_ready = dataUnits_44_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_45_ctrl_serveStealReq_ready = ctrlunits_45_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_45_ctrl_stealReq_ready = ctrlunits_45_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_45_data_availableTask_valid = dataUnits_45_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_45_data_availableTask_bits = dataUnits_45_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_45_data_qOutTask_ready = dataUnits_45_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_46_ctrl_serveStealReq_ready = ctrlunits_46_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_46_ctrl_stealReq_ready = ctrlunits_46_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_46_data_availableTask_valid = dataUnits_46_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_46_data_availableTask_bits = dataUnits_46_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_46_data_qOutTask_ready = dataUnits_46_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_47_ctrl_serveStealReq_ready = ctrlunits_47_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_47_ctrl_stealReq_ready = ctrlunits_47_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_47_data_availableTask_valid = dataUnits_47_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_47_data_availableTask_bits = dataUnits_47_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_47_data_qOutTask_ready = dataUnits_47_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_48_ctrl_serveStealReq_ready = ctrlunits_48_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_48_ctrl_stealReq_ready = ctrlunits_48_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_48_data_availableTask_valid = dataUnits_48_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_48_data_availableTask_bits = dataUnits_48_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_48_data_qOutTask_ready = dataUnits_48_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_49_ctrl_serveStealReq_ready = ctrlunits_49_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_49_ctrl_stealReq_ready = ctrlunits_49_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_49_data_availableTask_valid = dataUnits_49_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_49_data_availableTask_bits = dataUnits_49_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_49_data_qOutTask_ready = dataUnits_49_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_50_ctrl_serveStealReq_ready = ctrlunits_50_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_50_ctrl_stealReq_ready = ctrlunits_50_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_50_data_availableTask_valid = dataUnits_50_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_50_data_availableTask_bits = dataUnits_50_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_50_data_qOutTask_ready = dataUnits_50_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_51_ctrl_serveStealReq_ready = ctrlunits_51_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_51_ctrl_stealReq_ready = ctrlunits_51_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_51_data_availableTask_valid = dataUnits_51_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_51_data_availableTask_bits = dataUnits_51_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_51_data_qOutTask_ready = dataUnits_51_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_52_ctrl_serveStealReq_ready = ctrlunits_52_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_52_ctrl_stealReq_ready = ctrlunits_52_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_52_data_availableTask_valid = dataUnits_52_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_52_data_availableTask_bits = dataUnits_52_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_52_data_qOutTask_ready = dataUnits_52_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_53_ctrl_serveStealReq_ready = ctrlunits_53_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_53_ctrl_stealReq_ready = ctrlunits_53_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_53_data_availableTask_valid = dataUnits_53_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_53_data_availableTask_bits = dataUnits_53_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_53_data_qOutTask_ready = dataUnits_53_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_54_ctrl_serveStealReq_ready = ctrlunits_54_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_54_ctrl_stealReq_ready = ctrlunits_54_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_54_data_availableTask_valid = dataUnits_54_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_54_data_availableTask_bits = dataUnits_54_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_54_data_qOutTask_ready = dataUnits_54_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_55_ctrl_serveStealReq_ready = ctrlunits_55_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_55_ctrl_stealReq_ready = ctrlunits_55_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_55_data_availableTask_valid = dataUnits_55_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_55_data_availableTask_bits = dataUnits_55_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_55_data_qOutTask_ready = dataUnits_55_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_56_ctrl_serveStealReq_ready = ctrlunits_56_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_56_ctrl_stealReq_ready = ctrlunits_56_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_56_data_availableTask_valid = dataUnits_56_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_56_data_availableTask_bits = dataUnits_56_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_56_data_qOutTask_ready = dataUnits_56_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_57_ctrl_serveStealReq_ready = ctrlunits_57_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_57_ctrl_stealReq_ready = ctrlunits_57_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_57_data_availableTask_valid = dataUnits_57_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_57_data_availableTask_bits = dataUnits_57_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_57_data_qOutTask_ready = dataUnits_57_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_58_ctrl_serveStealReq_ready = ctrlunits_58_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_58_ctrl_stealReq_ready = ctrlunits_58_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_58_data_availableTask_valid = dataUnits_58_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_58_data_availableTask_bits = dataUnits_58_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_58_data_qOutTask_ready = dataUnits_58_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_59_ctrl_serveStealReq_ready = ctrlunits_59_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_59_ctrl_stealReq_ready = ctrlunits_59_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_59_data_availableTask_valid = dataUnits_59_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_59_data_availableTask_bits = dataUnits_59_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_59_data_qOutTask_ready = dataUnits_59_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_60_ctrl_serveStealReq_ready = ctrlunits_60_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_60_ctrl_stealReq_ready = ctrlunits_60_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_60_data_availableTask_valid = dataUnits_60_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_60_data_availableTask_bits = dataUnits_60_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_60_data_qOutTask_ready = dataUnits_60_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_61_ctrl_serveStealReq_ready = ctrlunits_61_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_61_ctrl_stealReq_ready = ctrlunits_61_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_61_data_availableTask_valid = dataUnits_61_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_61_data_availableTask_bits = dataUnits_61_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_61_data_qOutTask_ready = dataUnits_61_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_62_ctrl_serveStealReq_ready = ctrlunits_62_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_62_ctrl_stealReq_ready = ctrlunits_62_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_62_data_availableTask_valid = dataUnits_62_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_62_data_availableTask_bits = dataUnits_62_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_62_data_qOutTask_ready = dataUnits_62_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_63_ctrl_serveStealReq_ready = ctrlunits_63_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_63_ctrl_stealReq_ready = ctrlunits_63_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_63_data_availableTask_valid = dataUnits_63_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_63_data_availableTask_bits = dataUnits_63_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_63_data_qOutTask_ready = dataUnits_63_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_64_ctrl_serveStealReq_ready = ctrlunits_64_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_64_ctrl_stealReq_ready = ctrlunits_64_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_64_data_availableTask_valid = dataUnits_64_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_64_data_availableTask_bits = dataUnits_64_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_64_data_qOutTask_ready = dataUnits_64_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_65_ctrl_serveStealReq_ready = ctrlunits_65_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_65_ctrl_stealReq_ready = ctrlunits_65_io_connSS_stealReq_ready; // @[stealNetwork.scala 41:32]
  assign io_connSS_65_data_availableTask_valid = dataUnits_65_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_65_data_availableTask_bits = dataUnits_65_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_65_data_qOutTask_ready = dataUnits_65_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_connSS_66_ctrl_serveStealReq_ready = ctrlunits_66_io_connSS_serveStealReq_ready; // @[stealNetwork.scala 45:36]
  assign io_connSS_66_ctrl_stealReq_ready = ctrlunits_66_io_connSS_stealReq_ready; // @[stealNetwork.scala 45:36]
  assign io_connSS_66_data_availableTask_valid = dataUnits_66_io_connSS_availableTask_valid; // @[stealNetwork.scala 31:32]
  assign io_connSS_66_data_availableTask_bits = dataUnits_66_io_connSS_availableTask_bits; // @[stealNetwork.scala 31:32]
  assign io_connSS_66_data_qOutTask_ready = dataUnits_66_io_connSS_qOutTask_ready; // @[stealNetwork.scala 31:32]
  assign io_ntwDataUnitOccupancyVSS_0 = dataUnits_0_io_occupied; // @[stealNetwork.scala 49:54]
  assign dataUnits_0_clock = clock;
  assign dataUnits_0_reset = reset;
  assign dataUnits_0_io_taskIn = dataUnits_66_io_taskOut; // @[stealNetwork.scala 34:27]
  assign dataUnits_0_io_validIn = dataUnits_66_io_validOut; // @[stealNetwork.scala 35:27]
  assign dataUnits_0_io_connSS_availableTask_ready = io_connSS_0_data_availableTask_ready; // @[stealNetwork.scala 36:27]
  assign dataUnits_0_io_connSS_qOutTask_valid = io_connSS_0_data_qOutTask_valid; // @[stealNetwork.scala 36:27]
  assign dataUnits_0_io_connSS_qOutTask_bits = io_connSS_0_data_qOutTask_bits; // @[stealNetwork.scala 36:27]
  assign dataUnits_1_clock = clock;
  assign dataUnits_1_reset = reset;
  assign dataUnits_1_io_taskIn = dataUnits_0_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_1_io_validIn = dataUnits_0_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_1_io_connSS_availableTask_ready = 1'h0; // @[stealNetwork.scala 31:32]
  assign dataUnits_1_io_connSS_qOutTask_valid = io_connSS_1_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_1_io_connSS_qOutTask_bits = io_connSS_1_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_2_clock = clock;
  assign dataUnits_2_reset = reset;
  assign dataUnits_2_io_taskIn = dataUnits_1_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_2_io_validIn = dataUnits_1_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_2_io_connSS_availableTask_ready = 1'h0; // @[stealNetwork.scala 31:32]
  assign dataUnits_2_io_connSS_qOutTask_valid = io_connSS_2_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_2_io_connSS_qOutTask_bits = io_connSS_2_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_3_clock = clock;
  assign dataUnits_3_reset = reset;
  assign dataUnits_3_io_taskIn = dataUnits_2_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_3_io_validIn = dataUnits_2_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_3_io_connSS_availableTask_ready = io_connSS_3_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_3_io_connSS_qOutTask_valid = io_connSS_3_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_3_io_connSS_qOutTask_bits = io_connSS_3_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_4_clock = clock;
  assign dataUnits_4_reset = reset;
  assign dataUnits_4_io_taskIn = dataUnits_3_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_4_io_validIn = dataUnits_3_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_4_io_connSS_availableTask_ready = io_connSS_4_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_4_io_connSS_qOutTask_valid = io_connSS_4_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_4_io_connSS_qOutTask_bits = io_connSS_4_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_5_clock = clock;
  assign dataUnits_5_reset = reset;
  assign dataUnits_5_io_taskIn = dataUnits_4_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_5_io_validIn = dataUnits_4_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_5_io_connSS_availableTask_ready = io_connSS_5_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_5_io_connSS_qOutTask_valid = io_connSS_5_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_5_io_connSS_qOutTask_bits = io_connSS_5_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_6_clock = clock;
  assign dataUnits_6_reset = reset;
  assign dataUnits_6_io_taskIn = dataUnits_5_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_6_io_validIn = dataUnits_5_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_6_io_connSS_availableTask_ready = io_connSS_6_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_6_io_connSS_qOutTask_valid = io_connSS_6_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_6_io_connSS_qOutTask_bits = io_connSS_6_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_7_clock = clock;
  assign dataUnits_7_reset = reset;
  assign dataUnits_7_io_taskIn = dataUnits_6_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_7_io_validIn = dataUnits_6_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_7_io_connSS_availableTask_ready = io_connSS_7_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_7_io_connSS_qOutTask_valid = io_connSS_7_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_7_io_connSS_qOutTask_bits = io_connSS_7_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_8_clock = clock;
  assign dataUnits_8_reset = reset;
  assign dataUnits_8_io_taskIn = dataUnits_7_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_8_io_validIn = dataUnits_7_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_8_io_connSS_availableTask_ready = io_connSS_8_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_8_io_connSS_qOutTask_valid = io_connSS_8_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_8_io_connSS_qOutTask_bits = io_connSS_8_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_9_clock = clock;
  assign dataUnits_9_reset = reset;
  assign dataUnits_9_io_taskIn = dataUnits_8_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_9_io_validIn = dataUnits_8_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_9_io_connSS_availableTask_ready = io_connSS_9_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_9_io_connSS_qOutTask_valid = io_connSS_9_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_9_io_connSS_qOutTask_bits = io_connSS_9_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_10_clock = clock;
  assign dataUnits_10_reset = reset;
  assign dataUnits_10_io_taskIn = dataUnits_9_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_10_io_validIn = dataUnits_9_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_10_io_connSS_availableTask_ready = io_connSS_10_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_10_io_connSS_qOutTask_valid = io_connSS_10_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_10_io_connSS_qOutTask_bits = io_connSS_10_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_11_clock = clock;
  assign dataUnits_11_reset = reset;
  assign dataUnits_11_io_taskIn = dataUnits_10_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_11_io_validIn = dataUnits_10_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_11_io_connSS_availableTask_ready = io_connSS_11_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_11_io_connSS_qOutTask_valid = io_connSS_11_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_11_io_connSS_qOutTask_bits = io_connSS_11_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_12_clock = clock;
  assign dataUnits_12_reset = reset;
  assign dataUnits_12_io_taskIn = dataUnits_11_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_12_io_validIn = dataUnits_11_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_12_io_connSS_availableTask_ready = io_connSS_12_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_12_io_connSS_qOutTask_valid = io_connSS_12_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_12_io_connSS_qOutTask_bits = io_connSS_12_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_13_clock = clock;
  assign dataUnits_13_reset = reset;
  assign dataUnits_13_io_taskIn = dataUnits_12_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_13_io_validIn = dataUnits_12_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_13_io_connSS_availableTask_ready = io_connSS_13_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_13_io_connSS_qOutTask_valid = io_connSS_13_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_13_io_connSS_qOutTask_bits = io_connSS_13_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_14_clock = clock;
  assign dataUnits_14_reset = reset;
  assign dataUnits_14_io_taskIn = dataUnits_13_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_14_io_validIn = dataUnits_13_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_14_io_connSS_availableTask_ready = io_connSS_14_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_14_io_connSS_qOutTask_valid = io_connSS_14_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_14_io_connSS_qOutTask_bits = io_connSS_14_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_15_clock = clock;
  assign dataUnits_15_reset = reset;
  assign dataUnits_15_io_taskIn = dataUnits_14_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_15_io_validIn = dataUnits_14_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_15_io_connSS_availableTask_ready = io_connSS_15_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_15_io_connSS_qOutTask_valid = io_connSS_15_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_15_io_connSS_qOutTask_bits = io_connSS_15_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_16_clock = clock;
  assign dataUnits_16_reset = reset;
  assign dataUnits_16_io_taskIn = dataUnits_15_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_16_io_validIn = dataUnits_15_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_16_io_connSS_availableTask_ready = io_connSS_16_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_16_io_connSS_qOutTask_valid = io_connSS_16_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_16_io_connSS_qOutTask_bits = io_connSS_16_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_17_clock = clock;
  assign dataUnits_17_reset = reset;
  assign dataUnits_17_io_taskIn = dataUnits_16_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_17_io_validIn = dataUnits_16_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_17_io_connSS_availableTask_ready = io_connSS_17_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_17_io_connSS_qOutTask_valid = io_connSS_17_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_17_io_connSS_qOutTask_bits = io_connSS_17_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_18_clock = clock;
  assign dataUnits_18_reset = reset;
  assign dataUnits_18_io_taskIn = dataUnits_17_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_18_io_validIn = dataUnits_17_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_18_io_connSS_availableTask_ready = io_connSS_18_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_18_io_connSS_qOutTask_valid = io_connSS_18_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_18_io_connSS_qOutTask_bits = io_connSS_18_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_19_clock = clock;
  assign dataUnits_19_reset = reset;
  assign dataUnits_19_io_taskIn = dataUnits_18_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_19_io_validIn = dataUnits_18_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_19_io_connSS_availableTask_ready = io_connSS_19_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_19_io_connSS_qOutTask_valid = io_connSS_19_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_19_io_connSS_qOutTask_bits = io_connSS_19_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_20_clock = clock;
  assign dataUnits_20_reset = reset;
  assign dataUnits_20_io_taskIn = dataUnits_19_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_20_io_validIn = dataUnits_19_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_20_io_connSS_availableTask_ready = io_connSS_20_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_20_io_connSS_qOutTask_valid = io_connSS_20_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_20_io_connSS_qOutTask_bits = io_connSS_20_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_21_clock = clock;
  assign dataUnits_21_reset = reset;
  assign dataUnits_21_io_taskIn = dataUnits_20_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_21_io_validIn = dataUnits_20_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_21_io_connSS_availableTask_ready = io_connSS_21_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_21_io_connSS_qOutTask_valid = io_connSS_21_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_21_io_connSS_qOutTask_bits = io_connSS_21_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_22_clock = clock;
  assign dataUnits_22_reset = reset;
  assign dataUnits_22_io_taskIn = dataUnits_21_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_22_io_validIn = dataUnits_21_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_22_io_connSS_availableTask_ready = io_connSS_22_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_22_io_connSS_qOutTask_valid = io_connSS_22_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_22_io_connSS_qOutTask_bits = io_connSS_22_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_23_clock = clock;
  assign dataUnits_23_reset = reset;
  assign dataUnits_23_io_taskIn = dataUnits_22_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_23_io_validIn = dataUnits_22_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_23_io_connSS_availableTask_ready = io_connSS_23_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_23_io_connSS_qOutTask_valid = io_connSS_23_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_23_io_connSS_qOutTask_bits = io_connSS_23_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_24_clock = clock;
  assign dataUnits_24_reset = reset;
  assign dataUnits_24_io_taskIn = dataUnits_23_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_24_io_validIn = dataUnits_23_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_24_io_connSS_availableTask_ready = io_connSS_24_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_24_io_connSS_qOutTask_valid = io_connSS_24_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_24_io_connSS_qOutTask_bits = io_connSS_24_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_25_clock = clock;
  assign dataUnits_25_reset = reset;
  assign dataUnits_25_io_taskIn = dataUnits_24_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_25_io_validIn = dataUnits_24_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_25_io_connSS_availableTask_ready = io_connSS_25_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_25_io_connSS_qOutTask_valid = io_connSS_25_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_25_io_connSS_qOutTask_bits = io_connSS_25_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_26_clock = clock;
  assign dataUnits_26_reset = reset;
  assign dataUnits_26_io_taskIn = dataUnits_25_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_26_io_validIn = dataUnits_25_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_26_io_connSS_availableTask_ready = io_connSS_26_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_26_io_connSS_qOutTask_valid = io_connSS_26_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_26_io_connSS_qOutTask_bits = io_connSS_26_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_27_clock = clock;
  assign dataUnits_27_reset = reset;
  assign dataUnits_27_io_taskIn = dataUnits_26_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_27_io_validIn = dataUnits_26_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_27_io_connSS_availableTask_ready = io_connSS_27_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_27_io_connSS_qOutTask_valid = io_connSS_27_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_27_io_connSS_qOutTask_bits = io_connSS_27_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_28_clock = clock;
  assign dataUnits_28_reset = reset;
  assign dataUnits_28_io_taskIn = dataUnits_27_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_28_io_validIn = dataUnits_27_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_28_io_connSS_availableTask_ready = io_connSS_28_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_28_io_connSS_qOutTask_valid = io_connSS_28_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_28_io_connSS_qOutTask_bits = io_connSS_28_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_29_clock = clock;
  assign dataUnits_29_reset = reset;
  assign dataUnits_29_io_taskIn = dataUnits_28_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_29_io_validIn = dataUnits_28_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_29_io_connSS_availableTask_ready = io_connSS_29_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_29_io_connSS_qOutTask_valid = io_connSS_29_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_29_io_connSS_qOutTask_bits = io_connSS_29_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_30_clock = clock;
  assign dataUnits_30_reset = reset;
  assign dataUnits_30_io_taskIn = dataUnits_29_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_30_io_validIn = dataUnits_29_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_30_io_connSS_availableTask_ready = io_connSS_30_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_30_io_connSS_qOutTask_valid = io_connSS_30_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_30_io_connSS_qOutTask_bits = io_connSS_30_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_31_clock = clock;
  assign dataUnits_31_reset = reset;
  assign dataUnits_31_io_taskIn = dataUnits_30_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_31_io_validIn = dataUnits_30_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_31_io_connSS_availableTask_ready = io_connSS_31_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_31_io_connSS_qOutTask_valid = io_connSS_31_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_31_io_connSS_qOutTask_bits = io_connSS_31_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_32_clock = clock;
  assign dataUnits_32_reset = reset;
  assign dataUnits_32_io_taskIn = dataUnits_31_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_32_io_validIn = dataUnits_31_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_32_io_connSS_availableTask_ready = io_connSS_32_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_32_io_connSS_qOutTask_valid = io_connSS_32_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_32_io_connSS_qOutTask_bits = io_connSS_32_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_33_clock = clock;
  assign dataUnits_33_reset = reset;
  assign dataUnits_33_io_taskIn = dataUnits_32_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_33_io_validIn = dataUnits_32_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_33_io_connSS_availableTask_ready = io_connSS_33_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_33_io_connSS_qOutTask_valid = io_connSS_33_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_33_io_connSS_qOutTask_bits = io_connSS_33_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_34_clock = clock;
  assign dataUnits_34_reset = reset;
  assign dataUnits_34_io_taskIn = dataUnits_33_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_34_io_validIn = dataUnits_33_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_34_io_connSS_availableTask_ready = io_connSS_34_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_34_io_connSS_qOutTask_valid = io_connSS_34_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_34_io_connSS_qOutTask_bits = io_connSS_34_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_35_clock = clock;
  assign dataUnits_35_reset = reset;
  assign dataUnits_35_io_taskIn = dataUnits_34_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_35_io_validIn = dataUnits_34_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_35_io_connSS_availableTask_ready = io_connSS_35_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_35_io_connSS_qOutTask_valid = io_connSS_35_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_35_io_connSS_qOutTask_bits = io_connSS_35_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_36_clock = clock;
  assign dataUnits_36_reset = reset;
  assign dataUnits_36_io_taskIn = dataUnits_35_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_36_io_validIn = dataUnits_35_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_36_io_connSS_availableTask_ready = io_connSS_36_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_36_io_connSS_qOutTask_valid = io_connSS_36_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_36_io_connSS_qOutTask_bits = io_connSS_36_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_37_clock = clock;
  assign dataUnits_37_reset = reset;
  assign dataUnits_37_io_taskIn = dataUnits_36_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_37_io_validIn = dataUnits_36_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_37_io_connSS_availableTask_ready = io_connSS_37_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_37_io_connSS_qOutTask_valid = io_connSS_37_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_37_io_connSS_qOutTask_bits = io_connSS_37_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_38_clock = clock;
  assign dataUnits_38_reset = reset;
  assign dataUnits_38_io_taskIn = dataUnits_37_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_38_io_validIn = dataUnits_37_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_38_io_connSS_availableTask_ready = io_connSS_38_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_38_io_connSS_qOutTask_valid = io_connSS_38_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_38_io_connSS_qOutTask_bits = io_connSS_38_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_39_clock = clock;
  assign dataUnits_39_reset = reset;
  assign dataUnits_39_io_taskIn = dataUnits_38_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_39_io_validIn = dataUnits_38_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_39_io_connSS_availableTask_ready = io_connSS_39_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_39_io_connSS_qOutTask_valid = io_connSS_39_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_39_io_connSS_qOutTask_bits = io_connSS_39_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_40_clock = clock;
  assign dataUnits_40_reset = reset;
  assign dataUnits_40_io_taskIn = dataUnits_39_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_40_io_validIn = dataUnits_39_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_40_io_connSS_availableTask_ready = io_connSS_40_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_40_io_connSS_qOutTask_valid = io_connSS_40_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_40_io_connSS_qOutTask_bits = io_connSS_40_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_41_clock = clock;
  assign dataUnits_41_reset = reset;
  assign dataUnits_41_io_taskIn = dataUnits_40_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_41_io_validIn = dataUnits_40_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_41_io_connSS_availableTask_ready = io_connSS_41_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_41_io_connSS_qOutTask_valid = io_connSS_41_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_41_io_connSS_qOutTask_bits = io_connSS_41_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_42_clock = clock;
  assign dataUnits_42_reset = reset;
  assign dataUnits_42_io_taskIn = dataUnits_41_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_42_io_validIn = dataUnits_41_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_42_io_connSS_availableTask_ready = io_connSS_42_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_42_io_connSS_qOutTask_valid = io_connSS_42_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_42_io_connSS_qOutTask_bits = io_connSS_42_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_43_clock = clock;
  assign dataUnits_43_reset = reset;
  assign dataUnits_43_io_taskIn = dataUnits_42_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_43_io_validIn = dataUnits_42_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_43_io_connSS_availableTask_ready = io_connSS_43_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_43_io_connSS_qOutTask_valid = io_connSS_43_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_43_io_connSS_qOutTask_bits = io_connSS_43_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_44_clock = clock;
  assign dataUnits_44_reset = reset;
  assign dataUnits_44_io_taskIn = dataUnits_43_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_44_io_validIn = dataUnits_43_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_44_io_connSS_availableTask_ready = io_connSS_44_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_44_io_connSS_qOutTask_valid = io_connSS_44_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_44_io_connSS_qOutTask_bits = io_connSS_44_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_45_clock = clock;
  assign dataUnits_45_reset = reset;
  assign dataUnits_45_io_taskIn = dataUnits_44_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_45_io_validIn = dataUnits_44_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_45_io_connSS_availableTask_ready = io_connSS_45_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_45_io_connSS_qOutTask_valid = io_connSS_45_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_45_io_connSS_qOutTask_bits = io_connSS_45_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_46_clock = clock;
  assign dataUnits_46_reset = reset;
  assign dataUnits_46_io_taskIn = dataUnits_45_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_46_io_validIn = dataUnits_45_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_46_io_connSS_availableTask_ready = io_connSS_46_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_46_io_connSS_qOutTask_valid = io_connSS_46_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_46_io_connSS_qOutTask_bits = io_connSS_46_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_47_clock = clock;
  assign dataUnits_47_reset = reset;
  assign dataUnits_47_io_taskIn = dataUnits_46_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_47_io_validIn = dataUnits_46_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_47_io_connSS_availableTask_ready = io_connSS_47_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_47_io_connSS_qOutTask_valid = io_connSS_47_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_47_io_connSS_qOutTask_bits = io_connSS_47_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_48_clock = clock;
  assign dataUnits_48_reset = reset;
  assign dataUnits_48_io_taskIn = dataUnits_47_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_48_io_validIn = dataUnits_47_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_48_io_connSS_availableTask_ready = io_connSS_48_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_48_io_connSS_qOutTask_valid = io_connSS_48_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_48_io_connSS_qOutTask_bits = io_connSS_48_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_49_clock = clock;
  assign dataUnits_49_reset = reset;
  assign dataUnits_49_io_taskIn = dataUnits_48_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_49_io_validIn = dataUnits_48_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_49_io_connSS_availableTask_ready = io_connSS_49_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_49_io_connSS_qOutTask_valid = io_connSS_49_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_49_io_connSS_qOutTask_bits = io_connSS_49_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_50_clock = clock;
  assign dataUnits_50_reset = reset;
  assign dataUnits_50_io_taskIn = dataUnits_49_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_50_io_validIn = dataUnits_49_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_50_io_connSS_availableTask_ready = io_connSS_50_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_50_io_connSS_qOutTask_valid = io_connSS_50_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_50_io_connSS_qOutTask_bits = io_connSS_50_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_51_clock = clock;
  assign dataUnits_51_reset = reset;
  assign dataUnits_51_io_taskIn = dataUnits_50_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_51_io_validIn = dataUnits_50_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_51_io_connSS_availableTask_ready = io_connSS_51_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_51_io_connSS_qOutTask_valid = io_connSS_51_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_51_io_connSS_qOutTask_bits = io_connSS_51_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_52_clock = clock;
  assign dataUnits_52_reset = reset;
  assign dataUnits_52_io_taskIn = dataUnits_51_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_52_io_validIn = dataUnits_51_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_52_io_connSS_availableTask_ready = io_connSS_52_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_52_io_connSS_qOutTask_valid = io_connSS_52_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_52_io_connSS_qOutTask_bits = io_connSS_52_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_53_clock = clock;
  assign dataUnits_53_reset = reset;
  assign dataUnits_53_io_taskIn = dataUnits_52_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_53_io_validIn = dataUnits_52_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_53_io_connSS_availableTask_ready = io_connSS_53_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_53_io_connSS_qOutTask_valid = io_connSS_53_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_53_io_connSS_qOutTask_bits = io_connSS_53_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_54_clock = clock;
  assign dataUnits_54_reset = reset;
  assign dataUnits_54_io_taskIn = dataUnits_53_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_54_io_validIn = dataUnits_53_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_54_io_connSS_availableTask_ready = io_connSS_54_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_54_io_connSS_qOutTask_valid = io_connSS_54_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_54_io_connSS_qOutTask_bits = io_connSS_54_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_55_clock = clock;
  assign dataUnits_55_reset = reset;
  assign dataUnits_55_io_taskIn = dataUnits_54_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_55_io_validIn = dataUnits_54_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_55_io_connSS_availableTask_ready = io_connSS_55_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_55_io_connSS_qOutTask_valid = io_connSS_55_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_55_io_connSS_qOutTask_bits = io_connSS_55_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_56_clock = clock;
  assign dataUnits_56_reset = reset;
  assign dataUnits_56_io_taskIn = dataUnits_55_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_56_io_validIn = dataUnits_55_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_56_io_connSS_availableTask_ready = io_connSS_56_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_56_io_connSS_qOutTask_valid = io_connSS_56_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_56_io_connSS_qOutTask_bits = io_connSS_56_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_57_clock = clock;
  assign dataUnits_57_reset = reset;
  assign dataUnits_57_io_taskIn = dataUnits_56_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_57_io_validIn = dataUnits_56_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_57_io_connSS_availableTask_ready = io_connSS_57_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_57_io_connSS_qOutTask_valid = io_connSS_57_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_57_io_connSS_qOutTask_bits = io_connSS_57_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_58_clock = clock;
  assign dataUnits_58_reset = reset;
  assign dataUnits_58_io_taskIn = dataUnits_57_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_58_io_validIn = dataUnits_57_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_58_io_connSS_availableTask_ready = io_connSS_58_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_58_io_connSS_qOutTask_valid = io_connSS_58_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_58_io_connSS_qOutTask_bits = io_connSS_58_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_59_clock = clock;
  assign dataUnits_59_reset = reset;
  assign dataUnits_59_io_taskIn = dataUnits_58_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_59_io_validIn = dataUnits_58_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_59_io_connSS_availableTask_ready = io_connSS_59_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_59_io_connSS_qOutTask_valid = io_connSS_59_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_59_io_connSS_qOutTask_bits = io_connSS_59_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_60_clock = clock;
  assign dataUnits_60_reset = reset;
  assign dataUnits_60_io_taskIn = dataUnits_59_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_60_io_validIn = dataUnits_59_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_60_io_connSS_availableTask_ready = io_connSS_60_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_60_io_connSS_qOutTask_valid = io_connSS_60_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_60_io_connSS_qOutTask_bits = io_connSS_60_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_61_clock = clock;
  assign dataUnits_61_reset = reset;
  assign dataUnits_61_io_taskIn = dataUnits_60_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_61_io_validIn = dataUnits_60_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_61_io_connSS_availableTask_ready = io_connSS_61_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_61_io_connSS_qOutTask_valid = io_connSS_61_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_61_io_connSS_qOutTask_bits = io_connSS_61_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_62_clock = clock;
  assign dataUnits_62_reset = reset;
  assign dataUnits_62_io_taskIn = dataUnits_61_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_62_io_validIn = dataUnits_61_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_62_io_connSS_availableTask_ready = io_connSS_62_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_62_io_connSS_qOutTask_valid = io_connSS_62_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_62_io_connSS_qOutTask_bits = io_connSS_62_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_63_clock = clock;
  assign dataUnits_63_reset = reset;
  assign dataUnits_63_io_taskIn = dataUnits_62_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_63_io_validIn = dataUnits_62_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_63_io_connSS_availableTask_ready = io_connSS_63_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_63_io_connSS_qOutTask_valid = io_connSS_63_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_63_io_connSS_qOutTask_bits = io_connSS_63_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_64_clock = clock;
  assign dataUnits_64_reset = reset;
  assign dataUnits_64_io_taskIn = dataUnits_63_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_64_io_validIn = dataUnits_63_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_64_io_connSS_availableTask_ready = io_connSS_64_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_64_io_connSS_qOutTask_valid = io_connSS_64_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_64_io_connSS_qOutTask_bits = io_connSS_64_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_65_clock = clock;
  assign dataUnits_65_reset = reset;
  assign dataUnits_65_io_taskIn = dataUnits_64_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_65_io_validIn = dataUnits_64_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_65_io_connSS_availableTask_ready = io_connSS_65_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_65_io_connSS_qOutTask_valid = io_connSS_65_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_65_io_connSS_qOutTask_bits = io_connSS_65_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign dataUnits_66_clock = clock;
  assign dataUnits_66_reset = reset;
  assign dataUnits_66_io_taskIn = dataUnits_65_io_taskOut; // @[stealNetwork.scala 29:32]
  assign dataUnits_66_io_validIn = dataUnits_65_io_validOut; // @[stealNetwork.scala 30:32]
  assign dataUnits_66_io_connSS_availableTask_ready = io_connSS_66_data_availableTask_ready; // @[stealNetwork.scala 31:32]
  assign dataUnits_66_io_connSS_qOutTask_valid = io_connSS_66_data_qOutTask_valid; // @[stealNetwork.scala 31:32]
  assign dataUnits_66_io_connSS_qOutTask_bits = io_connSS_66_data_qOutTask_bits; // @[stealNetwork.scala 31:32]
  assign ctrlunits_0_clock = clock;
  assign ctrlunits_0_reset = reset;
  assign ctrlunits_0_io_reqTaskIn = ctrlunits_1_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_0_io_connSS_serveStealReq_valid = io_connSS_0_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_0_io_connSS_stealReq_valid = 1'h0; // @[stealNetwork.scala 41:32]
  assign ctrlunits_1_clock = clock;
  assign ctrlunits_1_reset = reset;
  assign ctrlunits_1_io_reqTaskIn = ctrlunits_2_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_1_io_connSS_serveStealReq_valid = io_connSS_1_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_1_io_connSS_stealReq_valid = 1'h0; // @[stealNetwork.scala 41:32]
  assign ctrlunits_2_clock = clock;
  assign ctrlunits_2_reset = reset;
  assign ctrlunits_2_io_reqTaskIn = ctrlunits_3_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_2_io_connSS_serveStealReq_valid = io_connSS_2_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_2_io_connSS_stealReq_valid = 1'h0; // @[stealNetwork.scala 41:32]
  assign ctrlunits_3_clock = clock;
  assign ctrlunits_3_reset = reset;
  assign ctrlunits_3_io_reqTaskIn = ctrlunits_4_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_3_io_connSS_serveStealReq_valid = io_connSS_3_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_3_io_connSS_stealReq_valid = io_connSS_3_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_4_clock = clock;
  assign ctrlunits_4_reset = reset;
  assign ctrlunits_4_io_reqTaskIn = ctrlunits_5_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_4_io_connSS_serveStealReq_valid = io_connSS_4_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_4_io_connSS_stealReq_valid = io_connSS_4_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_5_clock = clock;
  assign ctrlunits_5_reset = reset;
  assign ctrlunits_5_io_reqTaskIn = ctrlunits_6_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_5_io_connSS_serveStealReq_valid = io_connSS_5_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_5_io_connSS_stealReq_valid = io_connSS_5_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_6_clock = clock;
  assign ctrlunits_6_reset = reset;
  assign ctrlunits_6_io_reqTaskIn = ctrlunits_7_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_6_io_connSS_serveStealReq_valid = io_connSS_6_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_6_io_connSS_stealReq_valid = io_connSS_6_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_7_clock = clock;
  assign ctrlunits_7_reset = reset;
  assign ctrlunits_7_io_reqTaskIn = ctrlunits_8_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_7_io_connSS_serveStealReq_valid = io_connSS_7_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_7_io_connSS_stealReq_valid = io_connSS_7_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_8_clock = clock;
  assign ctrlunits_8_reset = reset;
  assign ctrlunits_8_io_reqTaskIn = ctrlunits_9_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_8_io_connSS_serveStealReq_valid = io_connSS_8_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_8_io_connSS_stealReq_valid = io_connSS_8_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_9_clock = clock;
  assign ctrlunits_9_reset = reset;
  assign ctrlunits_9_io_reqTaskIn = ctrlunits_10_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_9_io_connSS_serveStealReq_valid = io_connSS_9_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_9_io_connSS_stealReq_valid = io_connSS_9_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_10_clock = clock;
  assign ctrlunits_10_reset = reset;
  assign ctrlunits_10_io_reqTaskIn = ctrlunits_11_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_10_io_connSS_serveStealReq_valid = io_connSS_10_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_10_io_connSS_stealReq_valid = io_connSS_10_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_11_clock = clock;
  assign ctrlunits_11_reset = reset;
  assign ctrlunits_11_io_reqTaskIn = ctrlunits_12_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_11_io_connSS_serveStealReq_valid = io_connSS_11_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_11_io_connSS_stealReq_valid = io_connSS_11_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_12_clock = clock;
  assign ctrlunits_12_reset = reset;
  assign ctrlunits_12_io_reqTaskIn = ctrlunits_13_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_12_io_connSS_serveStealReq_valid = io_connSS_12_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_12_io_connSS_stealReq_valid = io_connSS_12_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_13_clock = clock;
  assign ctrlunits_13_reset = reset;
  assign ctrlunits_13_io_reqTaskIn = ctrlunits_14_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_13_io_connSS_serveStealReq_valid = io_connSS_13_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_13_io_connSS_stealReq_valid = io_connSS_13_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_14_clock = clock;
  assign ctrlunits_14_reset = reset;
  assign ctrlunits_14_io_reqTaskIn = ctrlunits_15_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_14_io_connSS_serveStealReq_valid = io_connSS_14_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_14_io_connSS_stealReq_valid = io_connSS_14_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_15_clock = clock;
  assign ctrlunits_15_reset = reset;
  assign ctrlunits_15_io_reqTaskIn = ctrlunits_16_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_15_io_connSS_serveStealReq_valid = io_connSS_15_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_15_io_connSS_stealReq_valid = io_connSS_15_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_16_clock = clock;
  assign ctrlunits_16_reset = reset;
  assign ctrlunits_16_io_reqTaskIn = ctrlunits_17_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_16_io_connSS_serveStealReq_valid = io_connSS_16_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_16_io_connSS_stealReq_valid = io_connSS_16_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_17_clock = clock;
  assign ctrlunits_17_reset = reset;
  assign ctrlunits_17_io_reqTaskIn = ctrlunits_18_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_17_io_connSS_serveStealReq_valid = io_connSS_17_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_17_io_connSS_stealReq_valid = io_connSS_17_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_18_clock = clock;
  assign ctrlunits_18_reset = reset;
  assign ctrlunits_18_io_reqTaskIn = ctrlunits_19_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_18_io_connSS_serveStealReq_valid = io_connSS_18_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_18_io_connSS_stealReq_valid = io_connSS_18_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_19_clock = clock;
  assign ctrlunits_19_reset = reset;
  assign ctrlunits_19_io_reqTaskIn = ctrlunits_20_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_19_io_connSS_serveStealReq_valid = io_connSS_19_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_19_io_connSS_stealReq_valid = io_connSS_19_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_20_clock = clock;
  assign ctrlunits_20_reset = reset;
  assign ctrlunits_20_io_reqTaskIn = ctrlunits_21_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_20_io_connSS_serveStealReq_valid = io_connSS_20_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_20_io_connSS_stealReq_valid = io_connSS_20_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_21_clock = clock;
  assign ctrlunits_21_reset = reset;
  assign ctrlunits_21_io_reqTaskIn = ctrlunits_22_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_21_io_connSS_serveStealReq_valid = io_connSS_21_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_21_io_connSS_stealReq_valid = io_connSS_21_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_22_clock = clock;
  assign ctrlunits_22_reset = reset;
  assign ctrlunits_22_io_reqTaskIn = ctrlunits_23_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_22_io_connSS_serveStealReq_valid = io_connSS_22_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_22_io_connSS_stealReq_valid = io_connSS_22_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_23_clock = clock;
  assign ctrlunits_23_reset = reset;
  assign ctrlunits_23_io_reqTaskIn = ctrlunits_24_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_23_io_connSS_serveStealReq_valid = io_connSS_23_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_23_io_connSS_stealReq_valid = io_connSS_23_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_24_clock = clock;
  assign ctrlunits_24_reset = reset;
  assign ctrlunits_24_io_reqTaskIn = ctrlunits_25_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_24_io_connSS_serveStealReq_valid = io_connSS_24_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_24_io_connSS_stealReq_valid = io_connSS_24_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_25_clock = clock;
  assign ctrlunits_25_reset = reset;
  assign ctrlunits_25_io_reqTaskIn = ctrlunits_26_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_25_io_connSS_serveStealReq_valid = io_connSS_25_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_25_io_connSS_stealReq_valid = io_connSS_25_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_26_clock = clock;
  assign ctrlunits_26_reset = reset;
  assign ctrlunits_26_io_reqTaskIn = ctrlunits_27_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_26_io_connSS_serveStealReq_valid = io_connSS_26_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_26_io_connSS_stealReq_valid = io_connSS_26_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_27_clock = clock;
  assign ctrlunits_27_reset = reset;
  assign ctrlunits_27_io_reqTaskIn = ctrlunits_28_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_27_io_connSS_serveStealReq_valid = io_connSS_27_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_27_io_connSS_stealReq_valid = io_connSS_27_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_28_clock = clock;
  assign ctrlunits_28_reset = reset;
  assign ctrlunits_28_io_reqTaskIn = ctrlunits_29_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_28_io_connSS_serveStealReq_valid = io_connSS_28_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_28_io_connSS_stealReq_valid = io_connSS_28_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_29_clock = clock;
  assign ctrlunits_29_reset = reset;
  assign ctrlunits_29_io_reqTaskIn = ctrlunits_30_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_29_io_connSS_serveStealReq_valid = io_connSS_29_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_29_io_connSS_stealReq_valid = io_connSS_29_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_30_clock = clock;
  assign ctrlunits_30_reset = reset;
  assign ctrlunits_30_io_reqTaskIn = ctrlunits_31_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_30_io_connSS_serveStealReq_valid = io_connSS_30_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_30_io_connSS_stealReq_valid = io_connSS_30_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_31_clock = clock;
  assign ctrlunits_31_reset = reset;
  assign ctrlunits_31_io_reqTaskIn = ctrlunits_32_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_31_io_connSS_serveStealReq_valid = io_connSS_31_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_31_io_connSS_stealReq_valid = io_connSS_31_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_32_clock = clock;
  assign ctrlunits_32_reset = reset;
  assign ctrlunits_32_io_reqTaskIn = ctrlunits_33_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_32_io_connSS_serveStealReq_valid = io_connSS_32_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_32_io_connSS_stealReq_valid = io_connSS_32_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_33_clock = clock;
  assign ctrlunits_33_reset = reset;
  assign ctrlunits_33_io_reqTaskIn = ctrlunits_34_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_33_io_connSS_serveStealReq_valid = io_connSS_33_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_33_io_connSS_stealReq_valid = io_connSS_33_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_34_clock = clock;
  assign ctrlunits_34_reset = reset;
  assign ctrlunits_34_io_reqTaskIn = ctrlunits_35_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_34_io_connSS_serveStealReq_valid = io_connSS_34_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_34_io_connSS_stealReq_valid = io_connSS_34_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_35_clock = clock;
  assign ctrlunits_35_reset = reset;
  assign ctrlunits_35_io_reqTaskIn = ctrlunits_36_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_35_io_connSS_serveStealReq_valid = io_connSS_35_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_35_io_connSS_stealReq_valid = io_connSS_35_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_36_clock = clock;
  assign ctrlunits_36_reset = reset;
  assign ctrlunits_36_io_reqTaskIn = ctrlunits_37_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_36_io_connSS_serveStealReq_valid = io_connSS_36_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_36_io_connSS_stealReq_valid = io_connSS_36_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_37_clock = clock;
  assign ctrlunits_37_reset = reset;
  assign ctrlunits_37_io_reqTaskIn = ctrlunits_38_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_37_io_connSS_serveStealReq_valid = io_connSS_37_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_37_io_connSS_stealReq_valid = io_connSS_37_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_38_clock = clock;
  assign ctrlunits_38_reset = reset;
  assign ctrlunits_38_io_reqTaskIn = ctrlunits_39_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_38_io_connSS_serveStealReq_valid = io_connSS_38_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_38_io_connSS_stealReq_valid = io_connSS_38_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_39_clock = clock;
  assign ctrlunits_39_reset = reset;
  assign ctrlunits_39_io_reqTaskIn = ctrlunits_40_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_39_io_connSS_serveStealReq_valid = io_connSS_39_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_39_io_connSS_stealReq_valid = io_connSS_39_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_40_clock = clock;
  assign ctrlunits_40_reset = reset;
  assign ctrlunits_40_io_reqTaskIn = ctrlunits_41_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_40_io_connSS_serveStealReq_valid = io_connSS_40_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_40_io_connSS_stealReq_valid = io_connSS_40_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_41_clock = clock;
  assign ctrlunits_41_reset = reset;
  assign ctrlunits_41_io_reqTaskIn = ctrlunits_42_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_41_io_connSS_serveStealReq_valid = io_connSS_41_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_41_io_connSS_stealReq_valid = io_connSS_41_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_42_clock = clock;
  assign ctrlunits_42_reset = reset;
  assign ctrlunits_42_io_reqTaskIn = ctrlunits_43_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_42_io_connSS_serveStealReq_valid = io_connSS_42_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_42_io_connSS_stealReq_valid = io_connSS_42_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_43_clock = clock;
  assign ctrlunits_43_reset = reset;
  assign ctrlunits_43_io_reqTaskIn = ctrlunits_44_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_43_io_connSS_serveStealReq_valid = io_connSS_43_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_43_io_connSS_stealReq_valid = io_connSS_43_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_44_clock = clock;
  assign ctrlunits_44_reset = reset;
  assign ctrlunits_44_io_reqTaskIn = ctrlunits_45_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_44_io_connSS_serveStealReq_valid = io_connSS_44_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_44_io_connSS_stealReq_valid = io_connSS_44_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_45_clock = clock;
  assign ctrlunits_45_reset = reset;
  assign ctrlunits_45_io_reqTaskIn = ctrlunits_46_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_45_io_connSS_serveStealReq_valid = io_connSS_45_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_45_io_connSS_stealReq_valid = io_connSS_45_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_46_clock = clock;
  assign ctrlunits_46_reset = reset;
  assign ctrlunits_46_io_reqTaskIn = ctrlunits_47_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_46_io_connSS_serveStealReq_valid = io_connSS_46_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_46_io_connSS_stealReq_valid = io_connSS_46_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_47_clock = clock;
  assign ctrlunits_47_reset = reset;
  assign ctrlunits_47_io_reqTaskIn = ctrlunits_48_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_47_io_connSS_serveStealReq_valid = io_connSS_47_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_47_io_connSS_stealReq_valid = io_connSS_47_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_48_clock = clock;
  assign ctrlunits_48_reset = reset;
  assign ctrlunits_48_io_reqTaskIn = ctrlunits_49_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_48_io_connSS_serveStealReq_valid = io_connSS_48_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_48_io_connSS_stealReq_valid = io_connSS_48_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_49_clock = clock;
  assign ctrlunits_49_reset = reset;
  assign ctrlunits_49_io_reqTaskIn = ctrlunits_50_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_49_io_connSS_serveStealReq_valid = io_connSS_49_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_49_io_connSS_stealReq_valid = io_connSS_49_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_50_clock = clock;
  assign ctrlunits_50_reset = reset;
  assign ctrlunits_50_io_reqTaskIn = ctrlunits_51_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_50_io_connSS_serveStealReq_valid = io_connSS_50_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_50_io_connSS_stealReq_valid = io_connSS_50_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_51_clock = clock;
  assign ctrlunits_51_reset = reset;
  assign ctrlunits_51_io_reqTaskIn = ctrlunits_52_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_51_io_connSS_serveStealReq_valid = io_connSS_51_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_51_io_connSS_stealReq_valid = io_connSS_51_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_52_clock = clock;
  assign ctrlunits_52_reset = reset;
  assign ctrlunits_52_io_reqTaskIn = ctrlunits_53_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_52_io_connSS_serveStealReq_valid = io_connSS_52_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_52_io_connSS_stealReq_valid = io_connSS_52_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_53_clock = clock;
  assign ctrlunits_53_reset = reset;
  assign ctrlunits_53_io_reqTaskIn = ctrlunits_54_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_53_io_connSS_serveStealReq_valid = io_connSS_53_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_53_io_connSS_stealReq_valid = io_connSS_53_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_54_clock = clock;
  assign ctrlunits_54_reset = reset;
  assign ctrlunits_54_io_reqTaskIn = ctrlunits_55_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_54_io_connSS_serveStealReq_valid = io_connSS_54_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_54_io_connSS_stealReq_valid = io_connSS_54_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_55_clock = clock;
  assign ctrlunits_55_reset = reset;
  assign ctrlunits_55_io_reqTaskIn = ctrlunits_56_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_55_io_connSS_serveStealReq_valid = io_connSS_55_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_55_io_connSS_stealReq_valid = io_connSS_55_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_56_clock = clock;
  assign ctrlunits_56_reset = reset;
  assign ctrlunits_56_io_reqTaskIn = ctrlunits_57_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_56_io_connSS_serveStealReq_valid = io_connSS_56_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_56_io_connSS_stealReq_valid = io_connSS_56_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_57_clock = clock;
  assign ctrlunits_57_reset = reset;
  assign ctrlunits_57_io_reqTaskIn = ctrlunits_58_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_57_io_connSS_serveStealReq_valid = io_connSS_57_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_57_io_connSS_stealReq_valid = io_connSS_57_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_58_clock = clock;
  assign ctrlunits_58_reset = reset;
  assign ctrlunits_58_io_reqTaskIn = ctrlunits_59_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_58_io_connSS_serveStealReq_valid = io_connSS_58_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_58_io_connSS_stealReq_valid = io_connSS_58_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_59_clock = clock;
  assign ctrlunits_59_reset = reset;
  assign ctrlunits_59_io_reqTaskIn = ctrlunits_60_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_59_io_connSS_serveStealReq_valid = io_connSS_59_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_59_io_connSS_stealReq_valid = io_connSS_59_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_60_clock = clock;
  assign ctrlunits_60_reset = reset;
  assign ctrlunits_60_io_reqTaskIn = ctrlunits_61_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_60_io_connSS_serveStealReq_valid = io_connSS_60_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_60_io_connSS_stealReq_valid = io_connSS_60_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_61_clock = clock;
  assign ctrlunits_61_reset = reset;
  assign ctrlunits_61_io_reqTaskIn = ctrlunits_62_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_61_io_connSS_serveStealReq_valid = io_connSS_61_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_61_io_connSS_stealReq_valid = io_connSS_61_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_62_clock = clock;
  assign ctrlunits_62_reset = reset;
  assign ctrlunits_62_io_reqTaskIn = ctrlunits_63_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_62_io_connSS_serveStealReq_valid = io_connSS_62_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_62_io_connSS_stealReq_valid = io_connSS_62_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_63_clock = clock;
  assign ctrlunits_63_reset = reset;
  assign ctrlunits_63_io_reqTaskIn = ctrlunits_64_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_63_io_connSS_serveStealReq_valid = io_connSS_63_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_63_io_connSS_stealReq_valid = io_connSS_63_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_64_clock = clock;
  assign ctrlunits_64_reset = reset;
  assign ctrlunits_64_io_reqTaskIn = ctrlunits_65_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_64_io_connSS_serveStealReq_valid = io_connSS_64_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_64_io_connSS_stealReq_valid = io_connSS_64_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_65_clock = clock;
  assign ctrlunits_65_reset = reset;
  assign ctrlunits_65_io_reqTaskIn = ctrlunits_66_io_reqTaskOut; // @[stealNetwork.scala 40:32]
  assign ctrlunits_65_io_connSS_serveStealReq_valid = io_connSS_65_ctrl_serveStealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_65_io_connSS_stealReq_valid = io_connSS_65_ctrl_stealReq_valid; // @[stealNetwork.scala 41:32]
  assign ctrlunits_66_clock = clock;
  assign ctrlunits_66_reset = reset;
  assign ctrlunits_66_io_reqTaskIn = ctrlunits_0_io_reqTaskOut; // @[stealNetwork.scala 44:36]
  assign ctrlunits_66_io_connSS_serveStealReq_valid = io_connSS_66_ctrl_serveStealReq_valid; // @[stealNetwork.scala 45:36]
  assign ctrlunits_66_io_connSS_stealReq_valid = io_connSS_66_ctrl_stealReq_valid; // @[stealNetwork.scala 45:36]
endmodule
module stealServer(
  input          clock,
  input          reset,
  input          io_connNetwork_ctrl_serveStealReq_ready,
  output         io_connNetwork_ctrl_serveStealReq_valid,
  input          io_connNetwork_ctrl_stealReq_ready,
  output         io_connNetwork_ctrl_stealReq_valid,
  output         io_connNetwork_data_availableTask_ready,
  input          io_connNetwork_data_availableTask_valid,
  input  [255:0] io_connNetwork_data_availableTask_bits,
  input          io_connNetwork_data_qOutTask_ready,
  output         io_connNetwork_data_qOutTask_valid,
  output [255:0] io_connNetwork_data_qOutTask_bits,
  input  [5:0]   io_connQ_currLength,
  input          io_connQ_push_ready,
  output         io_connQ_push_valid,
  output [255:0] io_connQ_push_bits,
  output         io_connQ_pop_ready,
  input          io_connQ_pop_valid,
  input  [255:0] io_connQ_pop_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [255:0] _RAND_1;
  reg [255:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] stateReg; // @[stealServer.scala 28:39]
  reg [255:0] stolenTaskReg; // @[stealServer.scala 29:39]
  reg [255:0] giveTaskReg; // @[stealServer.scala 30:39]
  reg [31:0] requestKilledCount; // @[stealServer.scala 37:37]
  reg [31:0] requestTaskCount; // @[stealServer.scala 52:35]
  wire  _T_1 = io_connQ_currLength < 6'h6; // @[stealServer.scala 57:42]
  wire [31:0] _requestTaskCount_T_1 = requestTaskCount + 32'h1; // @[stealServer.scala 61:75]
  wire  _T_2 = io_connQ_currLength > 6'h16; // @[stealServer.scala 62:48]
  wire [2:0] _GEN_0 = io_connQ_currLength > 6'h6 ? 3'h6 : 3'h0; // @[stealServer.scala 64:68 65:55 67:55]
  wire [31:0] _GEN_3 = io_connQ_currLength < 6'h6 ? 32'h45 : requestKilledCount; // @[stealServer.scala 37:37 57:62 59:55]
  wire [31:0] _GEN_5 = io_connQ_currLength < 6'h6 ? _requestTaskCount_T_1 : requestTaskCount; // @[stealServer.scala 52:35 57:62 61:55]
  wire  _T_4 = stateReg == 3'h2; // @[stealServer.scala 69:33]
  wire  _T_5 = io_connQ_currLength >= 6'h6; // @[stealServer.scala 74:48]
  wire  _T_6 = requestKilledCount == 32'h0; // @[stealServer.scala 76:47]
  wire [31:0] _GEN_6 = requestKilledCount == 32'h0 ? _requestTaskCount_T_1 : requestTaskCount; // @[stealServer.scala 52:35 76:55 77:58]
  wire [2:0] _GEN_7 = requestKilledCount == 32'h0 ? stateReg : 3'h2; // @[stealServer.scala 28:39 76:55 79:58]
  wire [2:0] _GEN_8 = io_connQ_currLength >= 6'h6 ? 3'h0 : _GEN_7; // @[stealServer.scala 74:69 75:55]
  wire [31:0] _GEN_9 = io_connQ_currLength >= 6'h6 ? requestTaskCount : _GEN_6; // @[stealServer.scala 52:35 74:69]
  wire [31:0] _GEN_12 = io_connNetwork_data_availableTask_valid ? requestTaskCount : _GEN_9; // @[stealServer.scala 52:35 71:62]
  wire [31:0] _requestKilledCount_T_3 = requestKilledCount - 32'h1; // @[stealServer.scala 83:80]
  wire  _T_8 = stateReg == 3'h3; // @[stealServer.scala 90:33]
  wire [2:0] _GEN_14 = io_connQ_currLength >= 6'h16 ? 3'h5 : 3'h3; // @[stealServer.scala 93:69 94:58 97:58]
  wire [255:0] _GEN_15 = io_connQ_currLength >= 6'h16 ? stolenTaskReg : giveTaskReg; // @[stealServer.scala 30:39 93:69 95:58]
  wire [2:0] _GEN_16 = io_connQ_push_ready ? 3'h0 : _GEN_14; // @[stealServer.scala 91:42 92:58]
  wire [255:0] _GEN_17 = io_connQ_push_ready ? giveTaskReg : _GEN_15; // @[stealServer.scala 30:39 91:42]
  wire  _T_10 = stateReg == 3'h4; // @[stealServer.scala 103:33]
  wire  _T_11 = io_connQ_currLength == 6'h0; // @[stealServer.scala 107:48]
  wire [2:0] _GEN_18 = io_connQ_currLength == 6'h0 ? 3'h2 : 3'h4; // @[stealServer.scala 107:56 108:58 112:58]
  wire [31:0] _GEN_19 = io_connQ_currLength == 6'h0 ? 32'h45 : requestKilledCount; // @[stealServer.scala 107:56 109:58 37:37]
  wire [31:0] _GEN_20 = io_connQ_currLength == 6'h0 ? _requestTaskCount_T_1 : requestTaskCount; // @[stealServer.scala 107:56 110:58 52:35]
  wire [2:0] _GEN_21 = io_connQ_pop_valid ? 3'h5 : _GEN_18; // @[stealServer.scala 104:41 105:58]
  wire [255:0] _GEN_22 = io_connQ_pop_valid ? io_connQ_pop_bits : giveTaskReg; // @[stealServer.scala 104:41 106:58 30:39]
  wire [31:0] _GEN_23 = io_connQ_pop_valid ? requestKilledCount : _GEN_19; // @[stealServer.scala 104:41 37:37]
  wire [31:0] _GEN_24 = io_connQ_pop_valid ? requestTaskCount : _GEN_20; // @[stealServer.scala 104:41 52:35]
  wire  _T_12 = stateReg == 3'h5; // @[stealServer.scala 117:33]
  wire [2:0] _GEN_26 = io_connNetwork_data_qOutTask_ready ? 3'h0 : 3'h5; // @[stealServer.scala 118:57 120:58 122:58]
  wire  _T_13 = stateReg == 3'h6; // @[stealServer.scala 128:33]
  wire  _T_16 = io_connNetwork_ctrl_serveStealReq_ready & _T_5; // @[stealServer.scala 130:58]
  wire  _T_17 = _T_2 | _T_16; // @[stealServer.scala 129:61]
  wire [31:0] _requestTaskCount_T_7 = requestTaskCount + 32'h2; // @[stealServer.scala 135:75]
  wire [2:0] _GEN_28 = _T_1 ? 3'h2 : 3'h6; // @[stealServer.scala 136:68 138:55 141:58]
  wire [31:0] _GEN_30 = _T_1 & io_connNetwork_ctrl_serveStealReq_ready ? 32'h45 : _GEN_3; // @[stealServer.scala 132:111 133:55]
  wire [2:0] _GEN_31 = _T_1 & io_connNetwork_ctrl_serveStealReq_ready ? 3'h2 : _GEN_28; // @[stealServer.scala 132:111 134:55]
  wire [31:0] _GEN_32 = _T_1 & io_connNetwork_ctrl_serveStealReq_ready ? _requestTaskCount_T_7 : _GEN_5; // @[stealServer.scala 132:111 135:55]
  wire [2:0] _GEN_33 = _T_17 ? 3'h4 : _GEN_31; // @[stealServer.scala 130:103 131:55]
  wire [31:0] _GEN_34 = _T_17 ? requestKilledCount : _GEN_30; // @[stealServer.scala 130:103 37:37]
  wire [31:0] _GEN_35 = _T_17 ? requestTaskCount : _GEN_32; // @[stealServer.scala 130:103 52:35]
  wire [2:0] _GEN_36 = stateReg == 3'h6 ? _GEN_33 : stateReg; // @[stealServer.scala 128:62 28:39]
  wire [31:0] _GEN_37 = stateReg == 3'h6 ? _GEN_34 : requestKilledCount; // @[stealServer.scala 128:62 37:37]
  wire [31:0] _GEN_38 = stateReg == 3'h6 ? _GEN_35 : requestTaskCount; // @[stealServer.scala 128:62 52:35]
  wire [2:0] _GEN_41 = stateReg == 3'h5 ? _GEN_26 : _GEN_36; // @[stealServer.scala 117:56]
  wire [255:0] _GEN_43 = stateReg == 3'h5 ? giveTaskReg : 256'h0; // @[stealServer.scala 117:56 126:59 47:47]
  wire [31:0] _GEN_44 = stateReg == 3'h5 ? requestKilledCount : _GEN_37; // @[stealServer.scala 117:56 37:37]
  wire [31:0] _GEN_45 = stateReg == 3'h5 ? requestTaskCount : _GEN_38; // @[stealServer.scala 117:56 52:35]
  wire  _GEN_46 = stateReg == 3'h5 ? 1'h0 : _T_13; // @[stealServer.scala 117:56 50:47]
  wire [2:0] _GEN_47 = stateReg == 3'h4 ? _GEN_21 : _GEN_41; // @[stealServer.scala 103:51]
  wire [255:0] _GEN_48 = stateReg == 3'h4 ? _GEN_22 : giveTaskReg; // @[stealServer.scala 103:51 30:39]
  wire [31:0] _GEN_49 = stateReg == 3'h4 ? _GEN_23 : _GEN_44; // @[stealServer.scala 103:51]
  wire [31:0] _GEN_50 = stateReg == 3'h4 ? _GEN_24 : _GEN_45; // @[stealServer.scala 103:51]
  wire  _GEN_53 = stateReg == 3'h4 ? 1'h0 : _T_12; // @[stealServer.scala 103:51 46:47]
  wire [255:0] _GEN_54 = stateReg == 3'h4 ? 256'h0 : _GEN_43; // @[stealServer.scala 103:51 47:47]
  wire  _GEN_55 = stateReg == 3'h4 ? 1'h0 : _GEN_46; // @[stealServer.scala 103:51 50:47]
  wire [255:0] _GEN_58 = stateReg == 3'h3 ? stolenTaskReg : 256'h0; // @[stealServer.scala 90:52 100:59 42:47]
  wire [31:0] _GEN_61 = stateReg == 3'h3 ? requestTaskCount : _GEN_50; // @[stealServer.scala 52:35 90:52]
  wire  _GEN_62 = stateReg == 3'h3 ? 1'h0 : _T_10; // @[stealServer.scala 41:47 90:52]
  wire  _GEN_64 = stateReg == 3'h3 ? 1'h0 : _GEN_53; // @[stealServer.scala 46:47 90:52]
  wire [255:0] _GEN_65 = stateReg == 3'h3 ? 256'h0 : _GEN_54; // @[stealServer.scala 47:47 90:52]
  wire  _GEN_66 = stateReg == 3'h3 ? 1'h0 : _GEN_55; // @[stealServer.scala 50:47 90:52]
  wire [31:0] _GEN_69 = stateReg == 3'h2 ? _GEN_12 : _GEN_61; // @[stealServer.scala 69:54]
  wire [255:0] _GEN_73 = stateReg == 3'h2 ? 256'h0 : _GEN_58; // @[stealServer.scala 42:47 69:54]
  wire  _GEN_74 = stateReg == 3'h2 ? 1'h0 : _T_8; // @[stealServer.scala 43:47 69:54]
  wire  _GEN_75 = stateReg == 3'h2 ? 1'h0 : _GEN_62; // @[stealServer.scala 41:47 69:54]
  wire  _GEN_77 = stateReg == 3'h2 ? 1'h0 : _GEN_64; // @[stealServer.scala 46:47 69:54]
  wire [255:0] _GEN_78 = stateReg == 3'h2 ? 256'h0 : _GEN_65; // @[stealServer.scala 47:47 69:54]
  wire  _GEN_79 = stateReg == 3'h2 ? 1'h0 : _GEN_66; // @[stealServer.scala 50:47 69:54]
  wire [31:0] _GEN_83 = stateReg == 3'h0 ? _GEN_5 : _GEN_69; // @[stealServer.scala 56:38]
  wire  _T_21 = requestTaskCount > 32'h0; // @[stealServer.scala 148:35]
  wire  _T_26 = _T_21 & ~(_T_13 & _T_1); // @[stealServer.scala 149:17]
  wire  _T_31 = _T_26 & ~(_T_10 & _T_11); // @[stealServer.scala 150:17]
  wire  _T_36 = _T_31 & ~(_T_4 & _T_6); // @[stealServer.scala 151:17]
  wire [31:0] _requestTaskCount_T_11 = requestTaskCount - 32'h1; // @[stealServer.scala 156:58]
  assign io_connNetwork_ctrl_serveStealReq_valid = stateReg == 3'h0 ? 1'h0 : _GEN_79; // @[stealServer.scala 56:38 50:47]
  assign io_connNetwork_ctrl_stealReq_valid = _T_31 & ~(_T_4 & _T_6); // @[stealServer.scala 151:17]
  assign io_connNetwork_data_availableTask_ready = stateReg == 3'h0 ? 1'h0 : _T_4; // @[stealServer.scala 56:38 45:47]
  assign io_connNetwork_data_qOutTask_valid = stateReg == 3'h0 ? 1'h0 : _GEN_77; // @[stealServer.scala 56:38 46:47]
  assign io_connNetwork_data_qOutTask_bits = stateReg == 3'h0 ? 256'h0 : _GEN_78; // @[stealServer.scala 56:38 47:47]
  assign io_connQ_push_valid = stateReg == 3'h0 ? 1'h0 : _GEN_74; // @[stealServer.scala 56:38 43:47]
  assign io_connQ_push_bits = stateReg == 3'h0 ? 256'h0 : _GEN_73; // @[stealServer.scala 56:38 42:47]
  assign io_connQ_pop_ready = stateReg == 3'h0 ? 1'h0 : _GEN_75; // @[stealServer.scala 56:38 41:47]
  always @(posedge clock) begin
    if (reset) begin // @[stealServer.scala 28:39]
      stateReg <= 3'h0; // @[stealServer.scala 28:39]
    end else if (stateReg == 3'h0) begin // @[stealServer.scala 56:38]
      if (io_connQ_currLength < 6'h6) begin // @[stealServer.scala 57:62]
        stateReg <= 3'h2; // @[stealServer.scala 60:55]
      end else if (io_connQ_currLength > 6'h16) begin // @[stealServer.scala 62:68]
        stateReg <= 3'h4; // @[stealServer.scala 63:55]
      end else begin
        stateReg <= _GEN_0;
      end
    end else if (stateReg == 3'h2) begin // @[stealServer.scala 69:54]
      if (io_connNetwork_data_availableTask_valid) begin // @[stealServer.scala 71:62]
        stateReg <= 3'h3; // @[stealServer.scala 72:58]
      end else begin
        stateReg <= _GEN_8;
      end
    end else if (stateReg == 3'h3) begin // @[stealServer.scala 90:52]
      stateReg <= _GEN_16;
    end else begin
      stateReg <= _GEN_47;
    end
    if (reset) begin // @[stealServer.scala 29:39]
      stolenTaskReg <= 256'h0; // @[stealServer.scala 29:39]
    end else if (!(stateReg == 3'h0)) begin // @[stealServer.scala 56:38]
      if (stateReg == 3'h2) begin // @[stealServer.scala 69:54]
        if (io_connNetwork_data_availableTask_valid) begin // @[stealServer.scala 71:62]
          stolenTaskReg <= io_connNetwork_data_availableTask_bits; // @[stealServer.scala 73:58]
        end
      end
    end
    if (reset) begin // @[stealServer.scala 30:39]
      giveTaskReg <= 256'h0; // @[stealServer.scala 30:39]
    end else if (!(stateReg == 3'h0)) begin // @[stealServer.scala 56:38]
      if (!(stateReg == 3'h2)) begin // @[stealServer.scala 69:54]
        if (stateReg == 3'h3) begin // @[stealServer.scala 90:52]
          giveTaskReg <= _GEN_17;
        end else begin
          giveTaskReg <= _GEN_48;
        end
      end
    end
    if (reset) begin // @[stealServer.scala 37:37]
      requestKilledCount <= 32'h43; // @[stealServer.scala 37:37]
    end else if (stateReg == 3'h0) begin // @[stealServer.scala 56:38]
      if (io_connQ_currLength < 6'h6) begin // @[stealServer.scala 57:62]
        requestKilledCount <= 32'h45; // @[stealServer.scala 59:55]
      end
    end else if (stateReg == 3'h2) begin // @[stealServer.scala 69:54]
      if (~io_connNetwork_ctrl_serveStealReq_ready) begin // @[stealServer.scala 82:63]
        requestKilledCount <= _requestKilledCount_T_3; // @[stealServer.scala 83:58]
      end else begin
        requestKilledCount <= 32'h45; // @[stealServer.scala 85:58]
      end
    end else if (!(stateReg == 3'h3)) begin // @[stealServer.scala 90:52]
      requestKilledCount <= _GEN_49;
    end
    if (reset) begin // @[stealServer.scala 52:35]
      requestTaskCount <= 32'h0; // @[stealServer.scala 52:35]
    end else if (_T_36) begin // @[stealServer.scala 153:13]
      if (io_connNetwork_ctrl_stealReq_ready) begin // @[stealServer.scala 155:57]
        requestTaskCount <= _requestTaskCount_T_11; // @[stealServer.scala 156:38]
      end else begin
        requestTaskCount <= _GEN_83;
      end
    end else begin
      requestTaskCount <= _GEN_83;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[2:0];
  _RAND_1 = {8{`RANDOM}};
  stolenTaskReg = _RAND_1[255:0];
  _RAND_2 = {8{`RANDOM}};
  giveTaskReg = _RAND_2[255:0];
  _RAND_3 = {1{`RANDOM}};
  requestKilledCount = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  requestTaskCount = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module hw_deque(
  input          clock,
  input          reset,
  output         io_connVec_0_push_ready,
  input          io_connVec_0_push_valid,
  input  [255:0] io_connVec_0_push_bits,
  input          io_connVec_0_pop_ready,
  output         io_connVec_0_pop_valid,
  output [255:0] io_connVec_0_pop_bits,
  output [6:0]   io_connVec_1_currLength,
  output         io_connVec_1_push_ready,
  input          io_connVec_1_push_valid,
  input  [255:0] io_connVec_1_push_bits,
  input          io_connVec_1_pop_ready,
  output         io_connVec_1_pop_valid,
  output [255:0] io_connVec_1_pop_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  bramMem_clk; // @[deque.scala 34:30]
  wire  bramMem_rst; // @[deque.scala 34:30]
  wire [8:0] bramMem_a_addr; // @[deque.scala 34:30]
  wire [255:0] bramMem_a_din; // @[deque.scala 34:30]
  wire  bramMem_a_wr; // @[deque.scala 34:30]
  wire [255:0] bramMem_a_dout; // @[deque.scala 34:30]
  wire [8:0] bramMem_b_addr; // @[deque.scala 34:30]
  wire [255:0] bramMem_b_din; // @[deque.scala 34:30]
  wire  bramMem_b_wr; // @[deque.scala 34:30]
  wire [255:0] bramMem_b_dout; // @[deque.scala 34:30]
  reg [6:0] sideReg_0; // @[deque.scala 23:35]
  reg [6:0] sideReg_1; // @[deque.scala 23:81]
  reg  readLatency_0; // @[deque.scala 29:43]
  reg  readLatency_1; // @[deque.scala 29:43]
  reg [1:0] writeLatency_0; // @[deque.scala 30:43]
  reg [1:0] writeLatency_1; // @[deque.scala 30:43]
  reg [2:0] stateRegs_0; // @[deque.scala 54:40]
  reg [2:0] stateRegs_1; // @[deque.scala 54:40]
  wire [6:0] _currLen_T_1 = 7'h22 + sideReg_1; // @[deque.scala 177:31]
  wire [6:0] _currLen_T_3 = _currLen_T_1 - sideReg_0; // @[deque.scala 177:44]
  wire [6:0] _currLen_T_5 = _currLen_T_3 - 7'h1; // @[deque.scala 177:58]
  wire [6:0] _currLen_T_7 = sideReg_1 - sideReg_0; // @[deque.scala 179:31]
  wire [6:0] _currLen_T_9 = _currLen_T_7 - 7'h1; // @[deque.scala 179:44]
  wire [6:0] currLen = sideReg_0 > sideReg_1 ? _currLen_T_5 : _currLen_T_9; // @[deque.scala 176:34 177:17 179:17]
  wire  _T_1 = currLen > 7'h1; // @[deque.scala 74:58]
  wire  _T_3 = stateRegs_1 == 3'h0; // @[deque.scala 74:109]
  wire  _T_5 = currLen > 7'h0; // @[deque.scala 74:135]
  wire  _T_9 = io_connVec_0_push_valid & currLen < 7'h22; // @[deque.scala 76:53]
  wire [1:0] _GEN_1 = io_connVec_0_pop_ready & currLen > 7'h1 | io_connVec_0_pop_ready & stateRegs_1 == 3'h0 & currLen
     > 7'h0 ? 2'h2 : {{1'd0}, _T_9}; // @[deque.scala 74:142 75:34]
  wire  _T_10 = stateRegs_0 == 3'h1; // @[deque.scala 93:33]
  wire [1:0] _writeLatency_0_T_1 = writeLatency_0 - 2'h1; // @[deque.scala 99:52]
  wire [1:0] _GEN_3 = writeLatency_0 == 2'h0 ? 2'h3 : 2'h1; // @[deque.scala 100:33 95:42 97:33]
  wire  _GEN_4 = ~readLatency_0 ? 1'h0 : readLatency_0 - 1'h1; // @[deque.scala 108:41 109:33 112:33]
  wire [2:0] _GEN_5 = ~readLatency_0 ? 3'h4 : 3'h2; // @[deque.scala 108:41 110:33 113:33]
  wire [6:0] _T_15 = 7'h22 - 7'h1; // @[deque.scala 118:48]
  wire [6:0] _bramMem_io_a_addr_T_1 = sideReg_0 + 7'h1; // @[deque.scala 121:54]
  wire [6:0] _GEN_6 = sideReg_0 == _T_15 ? 7'h0 : _bramMem_io_a_addr_T_1; // @[deque.scala 118:54 119:39 121:39]
  wire  _T_17 = stateRegs_0 == 3'h4; // @[deque.scala 130:33]
  wire  _T_21 = stateRegs_0 == 3'h3; // @[deque.scala 154:33]
  wire [6:0] _sideReg_0_T_5 = sideReg_0 - 7'h1; // @[deque.scala 163:46]
  wire [6:0] _GEN_9 = sideReg_0 == 7'h0 ? _T_15 : _sideReg_0_T_5; // @[deque.scala 160:41 161:32 163:32]
  wire [2:0] _GEN_10 = stateRegs_0 == 3'h3 ? 3'h0 : stateRegs_0; // @[deque.scala 154:48 156:38 54:40]
  wire [6:0] _GEN_11 = stateRegs_0 == 3'h3 ? _GEN_9 : sideReg_0; // @[deque.scala 154:48 23:35]
  wire [2:0] _GEN_13 = stateRegs_0 == 3'h4 ? 3'h0 : _GEN_10; // @[deque.scala 130:47 132:38]
  wire [6:0] _GEN_14 = stateRegs_0 == 3'h4 ? _GEN_6 : _GEN_11; // @[deque.scala 130:47]
  wire [27:0] _GEN_15 = stateRegs_0 == 3'h4 ? {{21'd0}, _GEN_6} : 28'hfffffff; // @[deque.scala 130:47 59:34]
  wire [255:0] _GEN_17 = stateRegs_0 == 3'h4 ? bramMem_a_dout : 256'h0; // @[deque.scala 130:47 153:38 67:34]
  wire  _GEN_18 = stateRegs_0 == 3'h4 ? 1'h0 : _T_21; // @[deque.scala 130:47 65:34]
  wire [27:0] _GEN_21 = stateRegs_0 == 3'h2 ? {{21'd0}, _GEN_6} : _GEN_15; // @[deque.scala 106:51]
  wire  _GEN_23 = stateRegs_0 == 3'h2 ? 1'h0 : _T_17; // @[deque.scala 106:51 66:34]
  wire [255:0] _GEN_24 = stateRegs_0 == 3'h2 ? 256'h0 : _GEN_17; // @[deque.scala 106:51 67:34]
  wire  _GEN_25 = stateRegs_0 == 3'h2 ? 1'h0 : _GEN_18; // @[deque.scala 106:51 65:34]
  wire [27:0] _GEN_28 = stateRegs_0 == 3'h1 ? {{21'd0}, sideReg_0} : _GEN_21; // @[deque.scala 103:38 93:52]
  wire  _GEN_32 = stateRegs_0 == 3'h1 ? 1'h0 : _GEN_23; // @[deque.scala 66:34 93:52]
  wire [255:0] _GEN_33 = stateRegs_0 == 3'h1 ? 256'h0 : _GEN_24; // @[deque.scala 67:34 93:52]
  wire  _GEN_34 = stateRegs_0 == 3'h1 ? 1'h0 : _GEN_25; // @[deque.scala 65:34 93:52]
  wire [27:0] _GEN_37 = stateRegs_0 == 3'h0 ? 28'hfffffff : _GEN_28; // @[deque.scala 59:34 71:42]
  wire [1:0] _GEN_44 = io_connVec_1_pop_ready & _T_1 | io_connVec_1_pop_ready & ~io_connVec_0_pop_ready & _T_5 &
    stateRegs_0 != 3'h4 ? 2'h2 : 2'h0; // @[deque.scala 84:175 88:34 90:34]
  wire [1:0] _GEN_45 = io_connVec_1_push_valid & currLen < _T_15 ? 2'h1 : _GEN_44; // @[deque.scala 82:79 83:34]
  wire  _T_37 = stateRegs_1 == 3'h1; // @[deque.scala 93:33]
  wire [1:0] _writeLatency_1_T_1 = writeLatency_1 - 2'h1; // @[deque.scala 99:52]
  wire [1:0] _GEN_47 = writeLatency_1 == 2'h0 ? 2'h3 : 2'h1; // @[deque.scala 100:33 95:42 97:33]
  wire  _GEN_48 = ~readLatency_1 ? 1'h0 : readLatency_1 - 1'h1; // @[deque.scala 108:41 109:33 112:33]
  wire [2:0] _GEN_49 = ~readLatency_1 ? 3'h4 : 3'h2; // @[deque.scala 108:41 110:33 113:33]
  wire [6:0] _bramMem_io_b_addr_T_3 = sideReg_1 - 7'h1; // @[deque.scala 127:54]
  wire [6:0] _GEN_50 = sideReg_1 == 7'h0 ? _T_15 : _bramMem_io_b_addr_T_3; // @[deque.scala 124:41 125:39 127:39]
  wire  _T_42 = stateRegs_1 == 3'h4; // @[deque.scala 130:33]
  wire  _T_44 = stateRegs_1 == 3'h3; // @[deque.scala 154:33]
  wire [6:0] _sideReg_1_T_5 = sideReg_1 + 7'h1; // @[deque.scala 169:46]
  wire [6:0] _GEN_53 = sideReg_1 == _T_15 ? 7'h0 : _sideReg_1_T_5; // @[deque.scala 166:56 167:32 169:32]
  wire [2:0] _GEN_54 = stateRegs_1 == 3'h3 ? 3'h0 : stateRegs_1; // @[deque.scala 154:48 156:38 54:40]
  wire [6:0] _GEN_55 = stateRegs_1 == 3'h3 ? _GEN_53 : sideReg_1; // @[deque.scala 154:48 23:81]
  wire [2:0] _GEN_57 = stateRegs_1 == 3'h4 ? 3'h0 : _GEN_54; // @[deque.scala 130:47 132:38]
  wire [6:0] _GEN_58 = stateRegs_1 == 3'h4 ? _GEN_50 : _GEN_55; // @[deque.scala 130:47]
  wire [27:0] _GEN_59 = stateRegs_1 == 3'h4 ? {{21'd0}, _GEN_50} : 28'hfffffff; // @[deque.scala 130:47 59:34]
  wire [255:0] _GEN_61 = stateRegs_1 == 3'h4 ? bramMem_b_dout : 256'h0; // @[deque.scala 130:47 153:38 67:34]
  wire  _GEN_62 = stateRegs_1 == 3'h4 ? 1'h0 : _T_44; // @[deque.scala 130:47 65:34]
  wire [27:0] _GEN_65 = stateRegs_1 == 3'h2 ? {{21'd0}, _GEN_50} : _GEN_59; // @[deque.scala 106:51]
  wire  _GEN_67 = stateRegs_1 == 3'h2 ? 1'h0 : _T_42; // @[deque.scala 106:51 66:34]
  wire [255:0] _GEN_68 = stateRegs_1 == 3'h2 ? 256'h0 : _GEN_61; // @[deque.scala 106:51 67:34]
  wire  _GEN_69 = stateRegs_1 == 3'h2 ? 1'h0 : _GEN_62; // @[deque.scala 106:51 65:34]
  wire [27:0] _GEN_72 = stateRegs_1 == 3'h1 ? {{21'd0}, sideReg_1} : _GEN_65; // @[deque.scala 103:38 93:52]
  wire  _GEN_76 = stateRegs_1 == 3'h1 ? 1'h0 : _GEN_67; // @[deque.scala 66:34 93:52]
  wire [255:0] _GEN_77 = stateRegs_1 == 3'h1 ? 256'h0 : _GEN_68; // @[deque.scala 67:34 93:52]
  wire  _GEN_78 = stateRegs_1 == 3'h1 ? 1'h0 : _GEN_69; // @[deque.scala 65:34 93:52]
  wire [27:0] _GEN_81 = _T_3 ? 28'hfffffff : _GEN_72; // @[deque.scala 59:34 71:42]
  DualPortBRAM #(.DATA(256), .ADDR(9)) bramMem ( // @[deque.scala 34:30]
    .clk(bramMem_clk),
    .rst(bramMem_rst),
    .a_addr(bramMem_a_addr),
    .a_din(bramMem_a_din),
    .a_wr(bramMem_a_wr),
    .a_dout(bramMem_a_dout),
    .b_addr(bramMem_b_addr),
    .b_din(bramMem_b_din),
    .b_wr(bramMem_b_wr),
    .b_dout(bramMem_b_dout)
  );
  assign io_connVec_0_push_ready = stateRegs_0 == 3'h0 ? 1'h0 : _GEN_34; // @[deque.scala 65:34 71:42]
  assign io_connVec_0_pop_valid = stateRegs_0 == 3'h0 ? 1'h0 : _GEN_32; // @[deque.scala 66:34 71:42]
  assign io_connVec_0_pop_bits = stateRegs_0 == 3'h0 ? 256'h0 : _GEN_33; // @[deque.scala 67:34 71:42]
  assign io_connVec_1_currLength = sideReg_0 > sideReg_1 ? _currLen_T_5 : _currLen_T_9; // @[deque.scala 176:34 177:17 179:17]
  assign io_connVec_1_push_ready = _T_3 ? 1'h0 : _GEN_78; // @[deque.scala 65:34 71:42]
  assign io_connVec_1_pop_valid = _T_3 ? 1'h0 : _GEN_76; // @[deque.scala 66:34 71:42]
  assign io_connVec_1_pop_bits = _T_3 ? 256'h0 : _GEN_77; // @[deque.scala 67:34 71:42]
  assign bramMem_clk = clock; // @[deque.scala 36:22]
  assign bramMem_rst = reset; // @[deque.scala 37:22]
  assign bramMem_a_addr = _GEN_37[8:0];
  assign bramMem_a_din = io_connVec_0_push_bits; // @[deque.scala 60:34]
  assign bramMem_a_wr = stateRegs_0 == 3'h0 ? 1'h0 : _T_10; // @[deque.scala 61:34 71:42]
  assign bramMem_b_addr = _GEN_81[8:0];
  assign bramMem_b_din = io_connVec_1_push_bits; // @[deque.scala 60:34]
  assign bramMem_b_wr = _T_3 ? 1'h0 : _T_37; // @[deque.scala 61:34 71:42]
  always @(posedge clock) begin
    if (reset) begin // @[deque.scala 23:35]
      sideReg_0 <= 7'h0; // @[deque.scala 23:35]
    end else if (!(stateRegs_0 == 3'h0)) begin // @[deque.scala 71:42]
      if (!(stateRegs_0 == 3'h1)) begin // @[deque.scala 93:52]
        if (!(stateRegs_0 == 3'h2)) begin // @[deque.scala 106:51]
          sideReg_0 <= _GEN_14;
        end
      end
    end
    if (reset) begin // @[deque.scala 23:81]
      sideReg_1 <= 7'h1; // @[deque.scala 23:81]
    end else if (!(_T_3)) begin // @[deque.scala 71:42]
      if (!(stateRegs_1 == 3'h1)) begin // @[deque.scala 93:52]
        if (!(stateRegs_1 == 3'h2)) begin // @[deque.scala 106:51]
          sideReg_1 <= _GEN_58;
        end
      end
    end
    if (reset) begin // @[deque.scala 29:43]
      readLatency_0 <= 1'h0; // @[deque.scala 29:43]
    end else if (!(stateRegs_0 == 3'h0)) begin // @[deque.scala 71:42]
      if (!(stateRegs_0 == 3'h1)) begin // @[deque.scala 93:52]
        if (stateRegs_0 == 3'h2) begin // @[deque.scala 106:51]
          readLatency_0 <= _GEN_4;
        end
      end
    end
    if (reset) begin // @[deque.scala 29:43]
      readLatency_1 <= 1'h0; // @[deque.scala 29:43]
    end else if (!(_T_3)) begin // @[deque.scala 71:42]
      if (!(stateRegs_1 == 3'h1)) begin // @[deque.scala 93:52]
        if (stateRegs_1 == 3'h2) begin // @[deque.scala 106:51]
          readLatency_1 <= _GEN_48;
        end
      end
    end
    if (reset) begin // @[deque.scala 30:43]
      writeLatency_0 <= 2'h1; // @[deque.scala 30:43]
    end else if (!(stateRegs_0 == 3'h0)) begin // @[deque.scala 71:42]
      if (stateRegs_0 == 3'h1) begin // @[deque.scala 93:52]
        if (writeLatency_0 == 2'h0) begin // @[deque.scala 95:42]
          writeLatency_0 <= 2'h1; // @[deque.scala 96:33]
        end else begin
          writeLatency_0 <= _writeLatency_0_T_1; // @[deque.scala 99:33]
        end
      end
    end
    if (reset) begin // @[deque.scala 30:43]
      writeLatency_1 <= 2'h1; // @[deque.scala 30:43]
    end else if (!(_T_3)) begin // @[deque.scala 71:42]
      if (stateRegs_1 == 3'h1) begin // @[deque.scala 93:52]
        if (writeLatency_1 == 2'h0) begin // @[deque.scala 95:42]
          writeLatency_1 <= 2'h1; // @[deque.scala 96:33]
        end else begin
          writeLatency_1 <= _writeLatency_1_T_1; // @[deque.scala 99:33]
        end
      end
    end
    if (reset) begin // @[deque.scala 54:40]
      stateRegs_0 <= 3'h0; // @[deque.scala 54:40]
    end else if (stateRegs_0 == 3'h0) begin // @[deque.scala 71:42]
      stateRegs_0 <= {{1'd0}, _GEN_1};
    end else if (stateRegs_0 == 3'h1) begin // @[deque.scala 93:52]
      stateRegs_0 <= {{1'd0}, _GEN_3};
    end else if (stateRegs_0 == 3'h2) begin // @[deque.scala 106:51]
      stateRegs_0 <= _GEN_5;
    end else begin
      stateRegs_0 <= _GEN_13;
    end
    if (reset) begin // @[deque.scala 54:40]
      stateRegs_1 <= 3'h0; // @[deque.scala 54:40]
    end else if (_T_3) begin // @[deque.scala 71:42]
      stateRegs_1 <= {{1'd0}, _GEN_45};
    end else if (stateRegs_1 == 3'h1) begin // @[deque.scala 93:52]
      stateRegs_1 <= {{1'd0}, _GEN_47};
    end else if (stateRegs_1 == 3'h2) begin // @[deque.scala 106:51]
      stateRegs_1 <= _GEN_49;
    end else begin
      stateRegs_1 <= _GEN_57;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sideReg_0 = _RAND_0[6:0];
  _RAND_1 = {1{`RANDOM}};
  sideReg_1 = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  readLatency_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  readLatency_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  writeLatency_0 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  writeLatency_1 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  stateRegs_0 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  stateRegs_1 = _RAND_7[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module stealNW_TQ(
  input          clock,
  input          reset,
  output         io_connPE_0_push_ready,
  input          io_connPE_0_push_valid,
  input  [255:0] io_connPE_0_push_bits,
  input          io_connPE_0_pop_ready,
  output         io_connPE_0_pop_valid,
  output [255:0] io_connPE_0_pop_bits,
  output         io_connPE_1_push_ready,
  input          io_connPE_1_push_valid,
  input  [255:0] io_connPE_1_push_bits,
  input          io_connPE_1_pop_ready,
  output         io_connPE_1_pop_valid,
  output [255:0] io_connPE_1_pop_bits,
  output         io_connPE_2_push_ready,
  input          io_connPE_2_push_valid,
  input  [255:0] io_connPE_2_push_bits,
  input          io_connPE_2_pop_ready,
  output         io_connPE_2_pop_valid,
  output [255:0] io_connPE_2_pop_bits,
  output         io_connPE_3_push_ready,
  input          io_connPE_3_push_valid,
  input  [255:0] io_connPE_3_push_bits,
  input          io_connPE_3_pop_ready,
  output         io_connPE_3_pop_valid,
  output [255:0] io_connPE_3_pop_bits,
  output         io_connPE_4_push_ready,
  input          io_connPE_4_push_valid,
  input  [255:0] io_connPE_4_push_bits,
  input          io_connPE_4_pop_ready,
  output         io_connPE_4_pop_valid,
  output [255:0] io_connPE_4_pop_bits,
  output         io_connPE_5_push_ready,
  input          io_connPE_5_push_valid,
  input  [255:0] io_connPE_5_push_bits,
  input          io_connPE_5_pop_ready,
  output         io_connPE_5_pop_valid,
  output [255:0] io_connPE_5_pop_bits,
  output         io_connPE_6_push_ready,
  input          io_connPE_6_push_valid,
  input  [255:0] io_connPE_6_push_bits,
  input          io_connPE_6_pop_ready,
  output         io_connPE_6_pop_valid,
  output [255:0] io_connPE_6_pop_bits,
  output         io_connPE_7_push_ready,
  input          io_connPE_7_push_valid,
  input  [255:0] io_connPE_7_push_bits,
  input          io_connPE_7_pop_ready,
  output         io_connPE_7_pop_valid,
  output [255:0] io_connPE_7_pop_bits,
  output         io_connPE_8_push_ready,
  input          io_connPE_8_push_valid,
  input  [255:0] io_connPE_8_push_bits,
  input          io_connPE_8_pop_ready,
  output         io_connPE_8_pop_valid,
  output [255:0] io_connPE_8_pop_bits,
  output         io_connPE_9_push_ready,
  input          io_connPE_9_push_valid,
  input  [255:0] io_connPE_9_push_bits,
  input          io_connPE_9_pop_ready,
  output         io_connPE_9_pop_valid,
  output [255:0] io_connPE_9_pop_bits,
  output         io_connPE_10_push_ready,
  input          io_connPE_10_push_valid,
  input  [255:0] io_connPE_10_push_bits,
  input          io_connPE_10_pop_ready,
  output         io_connPE_10_pop_valid,
  output [255:0] io_connPE_10_pop_bits,
  output         io_connPE_11_push_ready,
  input          io_connPE_11_push_valid,
  input  [255:0] io_connPE_11_push_bits,
  input          io_connPE_11_pop_ready,
  output         io_connPE_11_pop_valid,
  output [255:0] io_connPE_11_pop_bits,
  output         io_connPE_12_push_ready,
  input          io_connPE_12_push_valid,
  input  [255:0] io_connPE_12_push_bits,
  input          io_connPE_12_pop_ready,
  output         io_connPE_12_pop_valid,
  output [255:0] io_connPE_12_pop_bits,
  output         io_connPE_13_push_ready,
  input          io_connPE_13_push_valid,
  input  [255:0] io_connPE_13_push_bits,
  input          io_connPE_13_pop_ready,
  output         io_connPE_13_pop_valid,
  output [255:0] io_connPE_13_pop_bits,
  output         io_connPE_14_push_ready,
  input          io_connPE_14_push_valid,
  input  [255:0] io_connPE_14_push_bits,
  input          io_connPE_14_pop_ready,
  output         io_connPE_14_pop_valid,
  output [255:0] io_connPE_14_pop_bits,
  output         io_connPE_15_push_ready,
  input          io_connPE_15_push_valid,
  input  [255:0] io_connPE_15_push_bits,
  input          io_connPE_15_pop_ready,
  output         io_connPE_15_pop_valid,
  output [255:0] io_connPE_15_pop_bits,
  output         io_connPE_16_push_ready,
  input          io_connPE_16_push_valid,
  input  [255:0] io_connPE_16_push_bits,
  input          io_connPE_16_pop_ready,
  output         io_connPE_16_pop_valid,
  output [255:0] io_connPE_16_pop_bits,
  output         io_connPE_17_push_ready,
  input          io_connPE_17_push_valid,
  input  [255:0] io_connPE_17_push_bits,
  input          io_connPE_17_pop_ready,
  output         io_connPE_17_pop_valid,
  output [255:0] io_connPE_17_pop_bits,
  output         io_connPE_18_push_ready,
  input          io_connPE_18_push_valid,
  input  [255:0] io_connPE_18_push_bits,
  input          io_connPE_18_pop_ready,
  output         io_connPE_18_pop_valid,
  output [255:0] io_connPE_18_pop_bits,
  output         io_connPE_19_push_ready,
  input          io_connPE_19_push_valid,
  input  [255:0] io_connPE_19_push_bits,
  input          io_connPE_19_pop_ready,
  output         io_connPE_19_pop_valid,
  output [255:0] io_connPE_19_pop_bits,
  output         io_connPE_20_push_ready,
  input          io_connPE_20_push_valid,
  input  [255:0] io_connPE_20_push_bits,
  input          io_connPE_20_pop_ready,
  output         io_connPE_20_pop_valid,
  output [255:0] io_connPE_20_pop_bits,
  output         io_connPE_21_push_ready,
  input          io_connPE_21_push_valid,
  input  [255:0] io_connPE_21_push_bits,
  input          io_connPE_21_pop_ready,
  output         io_connPE_21_pop_valid,
  output [255:0] io_connPE_21_pop_bits,
  output         io_connPE_22_push_ready,
  input          io_connPE_22_push_valid,
  input  [255:0] io_connPE_22_push_bits,
  input          io_connPE_22_pop_ready,
  output         io_connPE_22_pop_valid,
  output [255:0] io_connPE_22_pop_bits,
  output         io_connPE_23_push_ready,
  input          io_connPE_23_push_valid,
  input  [255:0] io_connPE_23_push_bits,
  input          io_connPE_23_pop_ready,
  output         io_connPE_23_pop_valid,
  output [255:0] io_connPE_23_pop_bits,
  output         io_connPE_24_push_ready,
  input          io_connPE_24_push_valid,
  input  [255:0] io_connPE_24_push_bits,
  input          io_connPE_24_pop_ready,
  output         io_connPE_24_pop_valid,
  output [255:0] io_connPE_24_pop_bits,
  output         io_connPE_25_push_ready,
  input          io_connPE_25_push_valid,
  input  [255:0] io_connPE_25_push_bits,
  input          io_connPE_25_pop_ready,
  output         io_connPE_25_pop_valid,
  output [255:0] io_connPE_25_pop_bits,
  output         io_connPE_26_push_ready,
  input          io_connPE_26_push_valid,
  input  [255:0] io_connPE_26_push_bits,
  input          io_connPE_26_pop_ready,
  output         io_connPE_26_pop_valid,
  output [255:0] io_connPE_26_pop_bits,
  output         io_connPE_27_push_ready,
  input          io_connPE_27_push_valid,
  input  [255:0] io_connPE_27_push_bits,
  input          io_connPE_27_pop_ready,
  output         io_connPE_27_pop_valid,
  output [255:0] io_connPE_27_pop_bits,
  output         io_connPE_28_push_ready,
  input          io_connPE_28_push_valid,
  input  [255:0] io_connPE_28_push_bits,
  input          io_connPE_28_pop_ready,
  output         io_connPE_28_pop_valid,
  output [255:0] io_connPE_28_pop_bits,
  output         io_connPE_29_push_ready,
  input          io_connPE_29_push_valid,
  input  [255:0] io_connPE_29_push_bits,
  input          io_connPE_29_pop_ready,
  output         io_connPE_29_pop_valid,
  output [255:0] io_connPE_29_pop_bits,
  output         io_connPE_30_push_ready,
  input          io_connPE_30_push_valid,
  input  [255:0] io_connPE_30_push_bits,
  input          io_connPE_30_pop_ready,
  output         io_connPE_30_pop_valid,
  output [255:0] io_connPE_30_pop_bits,
  output         io_connPE_31_push_ready,
  input          io_connPE_31_push_valid,
  input  [255:0] io_connPE_31_push_bits,
  input          io_connPE_31_pop_ready,
  output         io_connPE_31_pop_valid,
  output [255:0] io_connPE_31_pop_bits,
  output         io_connPE_32_push_ready,
  input          io_connPE_32_push_valid,
  input  [255:0] io_connPE_32_push_bits,
  input          io_connPE_32_pop_ready,
  output         io_connPE_32_pop_valid,
  output [255:0] io_connPE_32_pop_bits,
  output         io_connPE_33_push_ready,
  input          io_connPE_33_push_valid,
  input  [255:0] io_connPE_33_push_bits,
  input          io_connPE_33_pop_ready,
  output         io_connPE_33_pop_valid,
  output [255:0] io_connPE_33_pop_bits,
  output         io_connPE_34_push_ready,
  input          io_connPE_34_push_valid,
  input  [255:0] io_connPE_34_push_bits,
  input          io_connPE_34_pop_ready,
  output         io_connPE_34_pop_valid,
  output [255:0] io_connPE_34_pop_bits,
  output         io_connPE_35_push_ready,
  input          io_connPE_35_push_valid,
  input  [255:0] io_connPE_35_push_bits,
  input          io_connPE_35_pop_ready,
  output         io_connPE_35_pop_valid,
  output [255:0] io_connPE_35_pop_bits,
  output         io_connPE_36_push_ready,
  input          io_connPE_36_push_valid,
  input  [255:0] io_connPE_36_push_bits,
  input          io_connPE_36_pop_ready,
  output         io_connPE_36_pop_valid,
  output [255:0] io_connPE_36_pop_bits,
  output         io_connPE_37_push_ready,
  input          io_connPE_37_push_valid,
  input  [255:0] io_connPE_37_push_bits,
  input          io_connPE_37_pop_ready,
  output         io_connPE_37_pop_valid,
  output [255:0] io_connPE_37_pop_bits,
  output         io_connPE_38_push_ready,
  input          io_connPE_38_push_valid,
  input  [255:0] io_connPE_38_push_bits,
  input          io_connPE_38_pop_ready,
  output         io_connPE_38_pop_valid,
  output [255:0] io_connPE_38_pop_bits,
  output         io_connPE_39_push_ready,
  input          io_connPE_39_push_valid,
  input  [255:0] io_connPE_39_push_bits,
  input          io_connPE_39_pop_ready,
  output         io_connPE_39_pop_valid,
  output [255:0] io_connPE_39_pop_bits,
  output         io_connPE_40_push_ready,
  input          io_connPE_40_push_valid,
  input  [255:0] io_connPE_40_push_bits,
  input          io_connPE_40_pop_ready,
  output         io_connPE_40_pop_valid,
  output [255:0] io_connPE_40_pop_bits,
  output         io_connPE_41_push_ready,
  input          io_connPE_41_push_valid,
  input  [255:0] io_connPE_41_push_bits,
  input          io_connPE_41_pop_ready,
  output         io_connPE_41_pop_valid,
  output [255:0] io_connPE_41_pop_bits,
  output         io_connPE_42_push_ready,
  input          io_connPE_42_push_valid,
  input  [255:0] io_connPE_42_push_bits,
  input          io_connPE_42_pop_ready,
  output         io_connPE_42_pop_valid,
  output [255:0] io_connPE_42_pop_bits,
  output         io_connPE_43_push_ready,
  input          io_connPE_43_push_valid,
  input  [255:0] io_connPE_43_push_bits,
  input          io_connPE_43_pop_ready,
  output         io_connPE_43_pop_valid,
  output [255:0] io_connPE_43_pop_bits,
  output         io_connPE_44_push_ready,
  input          io_connPE_44_push_valid,
  input  [255:0] io_connPE_44_push_bits,
  input          io_connPE_44_pop_ready,
  output         io_connPE_44_pop_valid,
  output [255:0] io_connPE_44_pop_bits,
  output         io_connPE_45_push_ready,
  input          io_connPE_45_push_valid,
  input  [255:0] io_connPE_45_push_bits,
  input          io_connPE_45_pop_ready,
  output         io_connPE_45_pop_valid,
  output [255:0] io_connPE_45_pop_bits,
  output         io_connPE_46_push_ready,
  input          io_connPE_46_push_valid,
  input  [255:0] io_connPE_46_push_bits,
  input          io_connPE_46_pop_ready,
  output         io_connPE_46_pop_valid,
  output [255:0] io_connPE_46_pop_bits,
  output         io_connPE_47_push_ready,
  input          io_connPE_47_push_valid,
  input  [255:0] io_connPE_47_push_bits,
  input          io_connPE_47_pop_ready,
  output         io_connPE_47_pop_valid,
  output [255:0] io_connPE_47_pop_bits,
  output         io_connPE_48_push_ready,
  input          io_connPE_48_push_valid,
  input  [255:0] io_connPE_48_push_bits,
  input          io_connPE_48_pop_ready,
  output         io_connPE_48_pop_valid,
  output [255:0] io_connPE_48_pop_bits,
  output         io_connPE_49_push_ready,
  input          io_connPE_49_push_valid,
  input  [255:0] io_connPE_49_push_bits,
  input          io_connPE_49_pop_ready,
  output         io_connPE_49_pop_valid,
  output [255:0] io_connPE_49_pop_bits,
  output         io_connPE_50_push_ready,
  input          io_connPE_50_push_valid,
  input  [255:0] io_connPE_50_push_bits,
  input          io_connPE_50_pop_ready,
  output         io_connPE_50_pop_valid,
  output [255:0] io_connPE_50_pop_bits,
  output         io_connPE_51_push_ready,
  input          io_connPE_51_push_valid,
  input  [255:0] io_connPE_51_push_bits,
  input          io_connPE_51_pop_ready,
  output         io_connPE_51_pop_valid,
  output [255:0] io_connPE_51_pop_bits,
  output         io_connPE_52_push_ready,
  input          io_connPE_52_push_valid,
  input  [255:0] io_connPE_52_push_bits,
  input          io_connPE_52_pop_ready,
  output         io_connPE_52_pop_valid,
  output [255:0] io_connPE_52_pop_bits,
  output         io_connPE_53_push_ready,
  input          io_connPE_53_push_valid,
  input  [255:0] io_connPE_53_push_bits,
  input          io_connPE_53_pop_ready,
  output         io_connPE_53_pop_valid,
  output [255:0] io_connPE_53_pop_bits,
  output         io_connPE_54_push_ready,
  input          io_connPE_54_push_valid,
  input  [255:0] io_connPE_54_push_bits,
  input          io_connPE_54_pop_ready,
  output         io_connPE_54_pop_valid,
  output [255:0] io_connPE_54_pop_bits,
  output         io_connPE_55_push_ready,
  input          io_connPE_55_push_valid,
  input  [255:0] io_connPE_55_push_bits,
  input          io_connPE_55_pop_ready,
  output         io_connPE_55_pop_valid,
  output [255:0] io_connPE_55_pop_bits,
  output         io_connPE_56_push_ready,
  input          io_connPE_56_push_valid,
  input  [255:0] io_connPE_56_push_bits,
  input          io_connPE_56_pop_ready,
  output         io_connPE_56_pop_valid,
  output [255:0] io_connPE_56_pop_bits,
  output         io_connPE_57_push_ready,
  input          io_connPE_57_push_valid,
  input  [255:0] io_connPE_57_push_bits,
  input          io_connPE_57_pop_ready,
  output         io_connPE_57_pop_valid,
  output [255:0] io_connPE_57_pop_bits,
  output         io_connPE_58_push_ready,
  input          io_connPE_58_push_valid,
  input  [255:0] io_connPE_58_push_bits,
  input          io_connPE_58_pop_ready,
  output         io_connPE_58_pop_valid,
  output [255:0] io_connPE_58_pop_bits,
  output         io_connPE_59_push_ready,
  input          io_connPE_59_push_valid,
  input  [255:0] io_connPE_59_push_bits,
  input          io_connPE_59_pop_ready,
  output         io_connPE_59_pop_valid,
  output [255:0] io_connPE_59_pop_bits,
  output         io_connPE_60_push_ready,
  input          io_connPE_60_push_valid,
  input  [255:0] io_connPE_60_push_bits,
  input          io_connPE_60_pop_ready,
  output         io_connPE_60_pop_valid,
  output [255:0] io_connPE_60_pop_bits,
  output         io_connPE_61_push_ready,
  input          io_connPE_61_push_valid,
  input  [255:0] io_connPE_61_push_bits,
  input          io_connPE_61_pop_ready,
  output         io_connPE_61_pop_valid,
  output [255:0] io_connPE_61_pop_bits,
  output         io_connPE_62_push_ready,
  input          io_connPE_62_push_valid,
  input  [255:0] io_connPE_62_push_bits,
  input          io_connPE_62_pop_ready,
  output         io_connPE_62_pop_valid,
  output [255:0] io_connPE_62_pop_bits,
  output         io_connPE_63_push_ready,
  input          io_connPE_63_push_valid,
  input  [255:0] io_connPE_63_push_bits,
  input          io_connPE_63_pop_ready,
  output         io_connPE_63_pop_valid,
  output [255:0] io_connPE_63_pop_bits,
  output         io_connVSS_0_ctrl_serveStealReq_ready,
  input          io_connVSS_0_ctrl_serveStealReq_valid,
  input          io_connVSS_0_data_availableTask_ready,
  output         io_connVSS_0_data_availableTask_valid,
  output [255:0] io_connVSS_0_data_availableTask_bits,
  output         io_connVSS_0_data_qOutTask_ready,
  input          io_connVSS_0_data_qOutTask_valid,
  input  [255:0] io_connVSS_0_data_qOutTask_bits,
  output         io_connVAS_0_ctrl_serveStealReq_ready,
  input          io_connVAS_0_ctrl_serveStealReq_valid,
  output         io_connVAS_0_data_qOutTask_ready,
  input          io_connVAS_0_data_qOutTask_valid,
  input  [255:0] io_connVAS_0_data_qOutTask_bits,
  output         io_connVAS_1_ctrl_serveStealReq_ready,
  input          io_connVAS_1_ctrl_serveStealReq_valid,
  output         io_connVAS_1_data_qOutTask_ready,
  input          io_connVAS_1_data_qOutTask_valid,
  input  [255:0] io_connVAS_1_data_qOutTask_bits,
  output         io_ntwDataUnitOccupancyVSS_0
);
  wire  stealNet_clock; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_reset; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_0_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_0_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_0_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_0_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_0_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_0_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_0_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_0_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_1_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_1_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_1_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_1_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_1_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_2_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_2_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_2_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_2_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_2_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_3_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_3_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_3_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_3_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_3_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_3_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_3_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_3_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_3_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_3_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_4_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_4_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_4_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_4_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_4_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_4_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_4_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_4_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_4_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_4_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_5_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_5_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_5_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_5_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_5_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_5_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_5_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_5_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_5_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_5_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_6_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_6_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_6_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_6_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_6_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_6_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_6_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_6_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_6_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_6_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_7_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_7_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_7_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_7_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_7_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_7_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_7_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_7_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_7_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_7_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_8_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_8_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_8_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_8_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_8_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_8_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_8_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_8_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_8_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_8_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_9_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_9_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_9_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_9_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_9_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_9_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_9_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_9_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_9_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_9_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_10_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_10_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_10_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_10_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_10_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_10_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_10_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_10_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_10_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_10_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_11_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_11_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_11_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_11_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_11_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_11_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_11_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_11_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_11_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_11_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_12_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_12_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_12_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_12_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_12_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_12_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_12_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_12_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_12_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_12_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_13_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_13_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_13_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_13_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_13_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_13_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_13_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_13_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_13_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_13_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_14_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_14_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_14_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_14_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_14_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_14_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_14_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_14_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_14_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_14_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_15_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_15_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_15_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_15_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_15_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_15_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_15_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_15_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_15_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_15_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_16_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_16_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_16_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_16_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_16_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_16_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_16_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_16_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_16_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_16_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_17_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_17_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_17_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_17_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_17_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_17_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_17_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_17_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_17_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_17_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_18_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_18_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_18_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_18_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_18_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_18_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_18_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_18_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_18_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_18_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_19_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_19_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_19_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_19_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_19_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_19_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_19_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_19_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_19_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_19_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_20_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_20_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_20_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_20_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_20_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_20_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_20_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_20_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_20_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_20_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_21_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_21_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_21_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_21_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_21_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_21_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_21_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_21_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_21_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_21_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_22_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_22_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_22_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_22_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_22_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_22_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_22_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_22_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_22_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_22_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_23_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_23_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_23_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_23_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_23_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_23_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_23_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_23_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_23_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_23_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_24_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_24_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_24_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_24_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_24_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_24_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_24_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_24_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_24_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_24_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_25_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_25_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_25_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_25_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_25_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_25_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_25_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_25_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_25_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_25_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_26_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_26_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_26_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_26_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_26_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_26_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_26_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_26_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_26_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_26_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_27_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_27_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_27_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_27_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_27_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_27_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_27_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_27_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_27_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_27_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_28_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_28_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_28_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_28_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_28_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_28_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_28_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_28_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_28_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_28_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_29_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_29_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_29_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_29_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_29_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_29_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_29_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_29_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_29_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_29_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_30_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_30_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_30_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_30_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_30_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_30_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_30_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_30_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_30_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_30_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_31_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_31_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_31_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_31_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_31_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_31_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_31_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_31_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_31_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_31_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_32_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_32_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_32_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_32_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_32_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_32_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_32_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_32_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_32_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_32_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_33_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_33_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_33_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_33_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_33_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_33_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_33_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_33_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_33_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_33_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_34_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_34_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_34_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_34_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_34_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_34_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_34_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_34_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_34_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_34_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_35_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_35_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_35_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_35_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_35_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_35_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_35_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_35_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_35_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_35_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_36_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_36_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_36_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_36_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_36_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_36_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_36_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_36_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_36_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_36_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_37_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_37_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_37_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_37_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_37_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_37_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_37_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_37_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_37_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_37_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_38_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_38_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_38_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_38_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_38_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_38_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_38_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_38_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_38_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_38_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_39_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_39_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_39_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_39_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_39_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_39_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_39_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_39_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_39_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_39_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_40_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_40_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_40_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_40_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_40_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_40_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_40_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_40_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_40_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_40_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_41_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_41_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_41_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_41_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_41_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_41_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_41_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_41_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_41_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_41_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_42_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_42_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_42_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_42_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_42_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_42_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_42_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_42_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_42_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_42_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_43_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_43_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_43_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_43_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_43_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_43_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_43_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_43_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_43_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_43_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_44_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_44_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_44_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_44_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_44_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_44_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_44_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_44_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_44_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_44_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_45_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_45_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_45_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_45_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_45_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_45_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_45_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_45_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_45_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_45_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_46_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_46_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_46_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_46_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_46_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_46_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_46_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_46_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_46_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_46_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_47_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_47_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_47_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_47_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_47_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_47_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_47_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_47_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_47_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_47_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_48_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_48_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_48_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_48_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_48_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_48_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_48_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_48_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_48_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_48_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_49_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_49_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_49_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_49_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_49_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_49_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_49_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_49_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_49_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_49_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_50_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_50_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_50_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_50_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_50_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_50_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_50_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_50_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_50_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_50_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_51_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_51_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_51_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_51_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_51_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_51_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_51_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_51_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_51_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_51_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_52_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_52_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_52_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_52_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_52_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_52_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_52_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_52_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_52_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_52_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_53_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_53_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_53_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_53_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_53_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_53_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_53_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_53_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_53_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_53_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_54_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_54_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_54_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_54_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_54_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_54_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_54_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_54_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_54_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_54_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_55_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_55_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_55_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_55_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_55_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_55_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_55_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_55_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_55_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_55_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_56_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_56_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_56_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_56_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_56_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_56_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_56_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_56_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_56_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_56_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_57_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_57_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_57_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_57_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_57_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_57_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_57_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_57_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_57_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_57_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_58_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_58_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_58_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_58_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_58_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_58_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_58_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_58_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_58_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_58_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_59_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_59_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_59_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_59_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_59_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_59_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_59_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_59_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_59_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_59_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_60_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_60_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_60_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_60_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_60_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_60_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_60_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_60_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_60_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_60_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_61_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_61_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_61_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_61_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_61_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_61_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_61_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_61_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_61_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_61_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_62_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_62_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_62_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_62_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_62_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_62_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_62_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_62_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_62_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_62_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_63_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_63_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_63_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_63_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_63_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_63_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_63_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_63_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_63_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_63_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_64_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_64_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_64_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_64_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_64_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_64_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_64_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_64_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_64_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_64_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_65_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_65_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_65_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_65_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_65_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_65_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_65_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_65_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_65_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_65_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_66_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_66_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_66_ctrl_stealReq_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_66_ctrl_stealReq_valid; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_66_data_availableTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_66_data_availableTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_66_data_availableTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_66_data_qOutTask_ready; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_connSS_66_data_qOutTask_valid; // @[stealNW_TQ.scala 36:30]
  wire [255:0] stealNet_io_connSS_66_data_qOutTask_bits; // @[stealNW_TQ.scala 36:30]
  wire  stealNet_io_ntwDataUnitOccupancyVSS_0; // @[stealNW_TQ.scala 36:30]
  wire  stealServers_0_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_0_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_0_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_0_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_0_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_0_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_0_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_0_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_0_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_0_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_0_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_0_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_0_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_0_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_0_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_0_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_0_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_0_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_0_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_1_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_1_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_1_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_1_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_1_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_1_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_1_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_1_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_1_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_1_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_1_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_1_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_1_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_1_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_1_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_1_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_1_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_1_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_1_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_2_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_2_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_2_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_2_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_2_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_2_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_2_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_2_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_2_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_2_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_2_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_2_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_2_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_2_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_2_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_2_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_2_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_2_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_2_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_3_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_3_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_3_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_3_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_3_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_3_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_3_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_3_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_3_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_3_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_3_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_3_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_3_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_3_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_3_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_3_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_3_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_3_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_3_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_4_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_4_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_4_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_4_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_4_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_4_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_4_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_4_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_4_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_4_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_4_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_4_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_4_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_4_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_4_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_4_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_4_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_4_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_4_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_5_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_5_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_5_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_5_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_5_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_5_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_5_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_5_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_5_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_5_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_5_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_5_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_5_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_5_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_5_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_5_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_5_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_5_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_5_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_6_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_6_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_6_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_6_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_6_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_6_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_6_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_6_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_6_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_6_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_6_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_6_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_6_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_6_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_6_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_6_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_6_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_6_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_6_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_7_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_7_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_7_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_7_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_7_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_7_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_7_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_7_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_7_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_7_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_7_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_7_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_7_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_7_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_7_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_7_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_7_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_7_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_7_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_8_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_8_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_8_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_8_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_8_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_8_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_8_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_8_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_8_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_8_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_8_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_8_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_8_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_8_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_8_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_8_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_8_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_8_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_8_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_9_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_9_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_9_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_9_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_9_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_9_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_9_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_9_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_9_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_9_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_9_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_9_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_9_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_9_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_9_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_9_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_9_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_9_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_9_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_10_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_10_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_10_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_10_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_10_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_10_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_10_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_10_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_10_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_10_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_10_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_10_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_10_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_10_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_10_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_10_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_10_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_10_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_10_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_11_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_11_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_11_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_11_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_11_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_11_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_11_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_11_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_11_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_11_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_11_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_11_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_11_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_11_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_11_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_11_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_11_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_11_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_11_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_12_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_12_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_12_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_12_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_12_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_12_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_12_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_12_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_12_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_12_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_12_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_12_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_12_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_12_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_12_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_12_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_12_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_12_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_12_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_13_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_13_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_13_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_13_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_13_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_13_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_13_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_13_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_13_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_13_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_13_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_13_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_13_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_13_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_13_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_13_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_13_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_13_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_13_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_14_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_14_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_14_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_14_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_14_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_14_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_14_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_14_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_14_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_14_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_14_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_14_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_14_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_14_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_14_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_14_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_14_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_14_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_14_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_15_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_15_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_15_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_15_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_15_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_15_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_15_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_15_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_15_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_15_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_15_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_15_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_15_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_15_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_15_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_15_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_15_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_15_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_15_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_16_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_16_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_16_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_16_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_16_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_16_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_16_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_16_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_16_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_16_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_16_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_16_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_16_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_16_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_16_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_16_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_16_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_16_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_16_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_17_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_17_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_17_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_17_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_17_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_17_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_17_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_17_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_17_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_17_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_17_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_17_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_17_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_17_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_17_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_17_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_17_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_17_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_17_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_18_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_18_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_18_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_18_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_18_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_18_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_18_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_18_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_18_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_18_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_18_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_18_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_18_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_18_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_18_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_18_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_18_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_18_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_18_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_19_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_19_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_19_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_19_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_19_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_19_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_19_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_19_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_19_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_19_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_19_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_19_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_19_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_19_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_19_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_19_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_19_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_19_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_19_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_20_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_20_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_20_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_20_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_20_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_20_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_20_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_20_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_20_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_20_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_20_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_20_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_20_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_20_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_20_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_20_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_20_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_20_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_20_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_21_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_21_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_21_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_21_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_21_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_21_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_21_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_21_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_21_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_21_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_21_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_21_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_21_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_21_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_21_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_21_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_21_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_21_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_21_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_22_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_22_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_22_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_22_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_22_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_22_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_22_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_22_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_22_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_22_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_22_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_22_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_22_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_22_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_22_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_22_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_22_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_22_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_22_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_23_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_23_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_23_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_23_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_23_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_23_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_23_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_23_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_23_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_23_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_23_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_23_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_23_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_23_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_23_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_23_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_23_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_23_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_23_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_24_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_24_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_24_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_24_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_24_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_24_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_24_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_24_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_24_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_24_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_24_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_24_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_24_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_24_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_24_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_24_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_24_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_24_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_24_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_25_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_25_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_25_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_25_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_25_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_25_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_25_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_25_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_25_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_25_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_25_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_25_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_25_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_25_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_25_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_25_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_25_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_25_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_25_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_26_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_26_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_26_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_26_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_26_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_26_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_26_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_26_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_26_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_26_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_26_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_26_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_26_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_26_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_26_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_26_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_26_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_26_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_26_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_27_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_27_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_27_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_27_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_27_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_27_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_27_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_27_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_27_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_27_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_27_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_27_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_27_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_27_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_27_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_27_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_27_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_27_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_27_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_28_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_28_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_28_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_28_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_28_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_28_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_28_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_28_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_28_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_28_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_28_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_28_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_28_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_28_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_28_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_28_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_28_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_28_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_28_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_29_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_29_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_29_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_29_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_29_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_29_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_29_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_29_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_29_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_29_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_29_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_29_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_29_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_29_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_29_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_29_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_29_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_29_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_29_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_30_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_30_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_30_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_30_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_30_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_30_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_30_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_30_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_30_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_30_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_30_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_30_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_30_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_30_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_30_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_30_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_30_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_30_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_30_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_31_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_31_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_31_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_31_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_31_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_31_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_31_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_31_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_31_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_31_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_31_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_31_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_31_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_31_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_31_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_31_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_31_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_31_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_31_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_32_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_32_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_32_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_32_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_32_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_32_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_32_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_32_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_32_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_32_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_32_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_32_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_32_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_32_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_32_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_32_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_32_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_32_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_32_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_33_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_33_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_33_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_33_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_33_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_33_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_33_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_33_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_33_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_33_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_33_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_33_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_33_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_33_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_33_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_33_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_33_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_33_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_33_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_34_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_34_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_34_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_34_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_34_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_34_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_34_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_34_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_34_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_34_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_34_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_34_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_34_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_34_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_34_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_34_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_34_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_34_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_34_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_35_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_35_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_35_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_35_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_35_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_35_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_35_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_35_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_35_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_35_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_35_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_35_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_35_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_35_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_35_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_35_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_35_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_35_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_35_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_36_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_36_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_36_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_36_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_36_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_36_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_36_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_36_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_36_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_36_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_36_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_36_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_36_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_36_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_36_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_36_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_36_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_36_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_36_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_37_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_37_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_37_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_37_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_37_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_37_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_37_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_37_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_37_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_37_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_37_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_37_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_37_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_37_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_37_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_37_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_37_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_37_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_37_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_38_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_38_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_38_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_38_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_38_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_38_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_38_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_38_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_38_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_38_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_38_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_38_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_38_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_38_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_38_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_38_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_38_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_38_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_38_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_39_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_39_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_39_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_39_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_39_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_39_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_39_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_39_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_39_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_39_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_39_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_39_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_39_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_39_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_39_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_39_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_39_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_39_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_39_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_40_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_40_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_40_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_40_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_40_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_40_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_40_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_40_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_40_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_40_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_40_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_40_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_40_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_40_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_40_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_40_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_40_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_40_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_40_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_41_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_41_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_41_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_41_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_41_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_41_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_41_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_41_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_41_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_41_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_41_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_41_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_41_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_41_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_41_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_41_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_41_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_41_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_41_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_42_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_42_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_42_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_42_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_42_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_42_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_42_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_42_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_42_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_42_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_42_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_42_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_42_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_42_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_42_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_42_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_42_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_42_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_42_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_43_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_43_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_43_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_43_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_43_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_43_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_43_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_43_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_43_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_43_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_43_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_43_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_43_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_43_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_43_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_43_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_43_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_43_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_43_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_44_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_44_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_44_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_44_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_44_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_44_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_44_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_44_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_44_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_44_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_44_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_44_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_44_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_44_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_44_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_44_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_44_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_44_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_44_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_45_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_45_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_45_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_45_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_45_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_45_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_45_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_45_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_45_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_45_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_45_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_45_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_45_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_45_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_45_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_45_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_45_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_45_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_45_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_46_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_46_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_46_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_46_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_46_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_46_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_46_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_46_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_46_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_46_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_46_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_46_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_46_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_46_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_46_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_46_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_46_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_46_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_46_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_47_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_47_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_47_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_47_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_47_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_47_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_47_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_47_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_47_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_47_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_47_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_47_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_47_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_47_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_47_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_47_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_47_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_47_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_47_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_48_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_48_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_48_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_48_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_48_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_48_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_48_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_48_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_48_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_48_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_48_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_48_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_48_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_48_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_48_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_48_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_48_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_48_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_48_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_49_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_49_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_49_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_49_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_49_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_49_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_49_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_49_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_49_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_49_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_49_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_49_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_49_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_49_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_49_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_49_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_49_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_49_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_49_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_50_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_50_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_50_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_50_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_50_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_50_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_50_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_50_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_50_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_50_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_50_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_50_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_50_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_50_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_50_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_50_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_50_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_50_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_50_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_51_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_51_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_51_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_51_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_51_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_51_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_51_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_51_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_51_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_51_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_51_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_51_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_51_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_51_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_51_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_51_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_51_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_51_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_51_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_52_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_52_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_52_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_52_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_52_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_52_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_52_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_52_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_52_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_52_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_52_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_52_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_52_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_52_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_52_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_52_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_52_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_52_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_52_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_53_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_53_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_53_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_53_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_53_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_53_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_53_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_53_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_53_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_53_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_53_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_53_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_53_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_53_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_53_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_53_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_53_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_53_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_53_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_54_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_54_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_54_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_54_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_54_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_54_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_54_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_54_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_54_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_54_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_54_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_54_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_54_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_54_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_54_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_54_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_54_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_54_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_54_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_55_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_55_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_55_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_55_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_55_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_55_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_55_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_55_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_55_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_55_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_55_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_55_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_55_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_55_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_55_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_55_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_55_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_55_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_55_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_56_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_56_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_56_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_56_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_56_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_56_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_56_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_56_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_56_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_56_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_56_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_56_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_56_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_56_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_56_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_56_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_56_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_56_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_56_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_57_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_57_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_57_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_57_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_57_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_57_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_57_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_57_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_57_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_57_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_57_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_57_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_57_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_57_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_57_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_57_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_57_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_57_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_57_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_58_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_58_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_58_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_58_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_58_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_58_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_58_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_58_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_58_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_58_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_58_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_58_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_58_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_58_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_58_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_58_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_58_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_58_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_58_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_59_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_59_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_59_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_59_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_59_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_59_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_59_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_59_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_59_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_59_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_59_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_59_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_59_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_59_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_59_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_59_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_59_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_59_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_59_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_60_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_60_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_60_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_60_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_60_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_60_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_60_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_60_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_60_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_60_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_60_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_60_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_60_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_60_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_60_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_60_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_60_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_60_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_60_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_61_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_61_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_61_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_61_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_61_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_61_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_61_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_61_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_61_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_61_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_61_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_61_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_61_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_61_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_61_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_61_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_61_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_61_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_61_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_62_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_62_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_62_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_62_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_62_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_62_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_62_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_62_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_62_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_62_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_62_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_62_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_62_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_62_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_62_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_62_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_62_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_62_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_62_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_63_clock; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_63_reset; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_63_io_connNetwork_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_63_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_63_io_connNetwork_ctrl_stealReq_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_63_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_63_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_63_io_connNetwork_data_availableTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_63_io_connNetwork_data_availableTask_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_63_io_connNetwork_data_qOutTask_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_63_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_63_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 54:49]
  wire [5:0] stealServers_63_io_connQ_currLength; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_63_io_connQ_push_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_63_io_connQ_push_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_63_io_connQ_push_bits; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_63_io_connQ_pop_ready; // @[stealNW_TQ.scala 54:49]
  wire  stealServers_63_io_connQ_pop_valid; // @[stealNW_TQ.scala 54:49]
  wire [255:0] stealServers_63_io_connQ_pop_bits; // @[stealNW_TQ.scala 54:49]
  wire  taskQueues_0_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_0_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_0_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_0_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_0_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_0_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_0_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_0_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_0_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_0_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_0_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_0_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_0_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_0_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_0_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_1_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_1_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_1_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_1_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_1_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_1_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_1_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_1_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_1_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_1_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_1_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_1_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_1_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_1_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_1_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_2_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_2_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_2_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_2_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_2_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_2_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_2_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_2_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_2_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_2_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_2_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_2_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_2_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_2_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_2_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_3_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_3_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_3_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_3_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_3_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_3_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_3_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_3_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_3_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_3_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_3_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_3_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_3_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_3_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_3_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_4_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_4_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_4_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_4_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_4_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_4_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_4_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_4_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_4_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_4_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_4_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_4_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_4_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_4_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_4_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_5_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_5_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_5_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_5_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_5_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_5_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_5_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_5_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_5_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_5_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_5_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_5_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_5_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_5_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_5_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_6_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_6_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_6_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_6_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_6_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_6_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_6_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_6_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_6_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_6_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_6_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_6_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_6_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_6_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_6_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_7_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_7_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_7_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_7_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_7_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_7_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_7_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_7_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_7_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_7_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_7_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_7_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_7_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_7_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_7_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_8_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_8_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_8_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_8_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_8_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_8_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_8_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_8_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_8_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_8_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_8_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_8_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_8_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_8_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_8_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_9_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_9_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_9_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_9_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_9_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_9_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_9_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_9_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_9_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_9_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_9_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_9_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_9_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_9_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_9_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_10_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_10_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_10_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_10_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_10_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_10_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_10_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_10_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_10_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_10_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_10_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_10_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_10_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_10_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_10_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_11_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_11_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_11_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_11_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_11_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_11_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_11_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_11_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_11_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_11_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_11_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_11_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_11_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_11_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_11_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_12_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_12_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_12_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_12_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_12_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_12_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_12_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_12_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_12_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_12_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_12_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_12_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_12_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_12_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_12_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_13_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_13_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_13_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_13_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_13_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_13_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_13_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_13_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_13_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_13_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_13_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_13_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_13_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_13_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_13_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_14_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_14_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_14_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_14_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_14_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_14_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_14_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_14_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_14_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_14_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_14_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_14_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_14_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_14_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_14_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_15_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_15_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_15_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_15_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_15_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_15_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_15_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_15_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_15_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_15_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_15_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_15_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_15_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_15_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_15_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_16_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_16_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_16_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_16_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_16_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_16_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_16_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_16_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_16_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_16_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_16_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_16_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_16_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_16_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_16_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_17_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_17_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_17_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_17_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_17_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_17_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_17_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_17_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_17_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_17_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_17_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_17_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_17_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_17_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_17_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_18_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_18_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_18_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_18_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_18_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_18_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_18_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_18_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_18_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_18_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_18_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_18_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_18_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_18_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_18_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_19_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_19_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_19_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_19_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_19_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_19_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_19_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_19_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_19_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_19_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_19_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_19_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_19_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_19_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_19_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_20_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_20_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_20_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_20_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_20_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_20_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_20_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_20_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_20_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_20_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_20_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_20_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_20_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_20_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_20_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_21_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_21_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_21_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_21_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_21_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_21_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_21_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_21_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_21_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_21_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_21_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_21_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_21_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_21_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_21_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_22_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_22_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_22_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_22_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_22_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_22_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_22_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_22_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_22_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_22_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_22_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_22_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_22_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_22_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_22_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_23_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_23_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_23_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_23_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_23_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_23_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_23_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_23_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_23_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_23_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_23_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_23_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_23_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_23_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_23_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_24_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_24_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_24_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_24_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_24_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_24_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_24_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_24_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_24_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_24_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_24_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_24_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_24_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_24_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_24_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_25_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_25_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_25_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_25_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_25_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_25_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_25_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_25_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_25_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_25_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_25_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_25_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_25_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_25_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_25_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_26_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_26_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_26_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_26_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_26_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_26_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_26_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_26_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_26_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_26_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_26_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_26_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_26_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_26_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_26_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_27_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_27_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_27_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_27_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_27_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_27_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_27_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_27_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_27_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_27_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_27_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_27_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_27_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_27_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_27_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_28_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_28_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_28_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_28_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_28_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_28_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_28_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_28_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_28_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_28_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_28_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_28_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_28_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_28_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_28_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_29_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_29_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_29_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_29_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_29_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_29_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_29_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_29_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_29_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_29_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_29_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_29_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_29_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_29_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_29_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_30_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_30_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_30_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_30_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_30_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_30_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_30_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_30_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_30_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_30_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_30_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_30_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_30_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_30_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_30_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_31_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_31_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_31_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_31_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_31_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_31_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_31_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_31_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_31_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_31_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_31_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_31_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_31_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_31_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_31_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_32_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_32_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_32_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_32_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_32_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_32_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_32_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_32_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_32_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_32_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_32_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_32_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_32_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_32_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_32_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_33_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_33_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_33_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_33_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_33_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_33_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_33_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_33_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_33_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_33_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_33_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_33_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_33_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_33_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_33_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_34_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_34_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_34_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_34_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_34_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_34_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_34_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_34_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_34_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_34_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_34_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_34_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_34_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_34_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_34_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_35_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_35_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_35_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_35_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_35_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_35_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_35_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_35_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_35_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_35_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_35_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_35_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_35_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_35_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_35_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_36_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_36_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_36_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_36_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_36_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_36_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_36_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_36_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_36_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_36_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_36_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_36_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_36_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_36_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_36_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_37_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_37_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_37_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_37_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_37_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_37_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_37_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_37_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_37_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_37_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_37_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_37_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_37_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_37_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_37_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_38_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_38_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_38_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_38_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_38_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_38_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_38_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_38_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_38_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_38_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_38_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_38_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_38_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_38_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_38_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_39_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_39_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_39_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_39_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_39_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_39_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_39_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_39_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_39_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_39_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_39_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_39_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_39_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_39_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_39_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_40_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_40_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_40_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_40_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_40_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_40_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_40_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_40_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_40_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_40_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_40_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_40_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_40_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_40_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_40_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_41_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_41_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_41_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_41_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_41_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_41_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_41_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_41_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_41_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_41_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_41_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_41_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_41_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_41_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_41_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_42_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_42_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_42_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_42_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_42_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_42_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_42_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_42_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_42_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_42_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_42_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_42_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_42_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_42_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_42_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_43_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_43_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_43_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_43_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_43_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_43_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_43_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_43_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_43_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_43_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_43_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_43_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_43_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_43_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_43_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_44_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_44_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_44_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_44_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_44_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_44_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_44_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_44_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_44_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_44_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_44_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_44_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_44_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_44_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_44_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_45_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_45_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_45_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_45_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_45_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_45_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_45_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_45_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_45_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_45_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_45_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_45_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_45_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_45_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_45_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_46_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_46_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_46_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_46_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_46_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_46_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_46_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_46_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_46_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_46_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_46_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_46_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_46_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_46_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_46_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_47_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_47_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_47_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_47_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_47_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_47_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_47_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_47_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_47_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_47_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_47_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_47_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_47_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_47_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_47_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_48_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_48_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_48_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_48_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_48_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_48_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_48_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_48_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_48_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_48_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_48_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_48_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_48_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_48_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_48_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_49_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_49_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_49_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_49_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_49_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_49_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_49_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_49_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_49_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_49_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_49_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_49_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_49_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_49_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_49_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_50_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_50_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_50_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_50_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_50_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_50_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_50_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_50_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_50_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_50_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_50_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_50_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_50_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_50_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_50_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_51_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_51_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_51_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_51_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_51_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_51_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_51_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_51_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_51_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_51_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_51_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_51_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_51_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_51_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_51_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_52_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_52_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_52_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_52_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_52_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_52_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_52_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_52_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_52_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_52_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_52_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_52_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_52_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_52_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_52_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_53_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_53_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_53_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_53_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_53_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_53_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_53_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_53_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_53_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_53_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_53_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_53_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_53_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_53_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_53_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_54_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_54_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_54_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_54_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_54_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_54_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_54_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_54_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_54_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_54_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_54_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_54_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_54_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_54_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_54_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_55_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_55_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_55_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_55_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_55_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_55_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_55_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_55_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_55_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_55_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_55_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_55_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_55_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_55_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_55_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_56_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_56_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_56_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_56_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_56_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_56_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_56_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_56_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_56_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_56_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_56_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_56_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_56_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_56_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_56_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_57_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_57_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_57_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_57_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_57_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_57_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_57_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_57_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_57_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_57_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_57_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_57_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_57_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_57_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_57_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_58_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_58_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_58_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_58_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_58_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_58_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_58_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_58_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_58_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_58_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_58_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_58_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_58_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_58_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_58_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_59_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_59_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_59_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_59_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_59_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_59_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_59_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_59_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_59_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_59_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_59_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_59_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_59_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_59_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_59_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_60_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_60_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_60_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_60_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_60_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_60_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_60_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_60_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_60_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_60_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_60_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_60_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_60_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_60_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_60_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_61_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_61_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_61_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_61_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_61_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_61_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_61_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_61_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_61_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_61_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_61_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_61_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_61_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_61_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_61_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_62_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_62_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_62_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_62_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_62_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_62_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_62_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_62_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_62_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_62_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_62_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_62_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_62_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_62_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_62_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_63_clock; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_63_reset; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_63_io_connVec_0_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_63_io_connVec_0_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_63_io_connVec_0_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_63_io_connVec_0_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_63_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_63_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 58:49]
  wire [6:0] taskQueues_63_io_connVec_1_currLength; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_63_io_connVec_1_push_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_63_io_connVec_1_push_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_63_io_connVec_1_push_bits; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_63_io_connVec_1_pop_ready; // @[stealNW_TQ.scala 58:49]
  wire  taskQueues_63_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 58:49]
  wire [255:0] taskQueues_63_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 58:49]
  stealNetwork stealNet ( // @[stealNW_TQ.scala 36:30]
    .clock(stealNet_clock),
    .reset(stealNet_reset),
    .io_connSS_0_ctrl_serveStealReq_ready(stealNet_io_connSS_0_ctrl_serveStealReq_ready),
    .io_connSS_0_ctrl_serveStealReq_valid(stealNet_io_connSS_0_ctrl_serveStealReq_valid),
    .io_connSS_0_data_availableTask_ready(stealNet_io_connSS_0_data_availableTask_ready),
    .io_connSS_0_data_availableTask_valid(stealNet_io_connSS_0_data_availableTask_valid),
    .io_connSS_0_data_availableTask_bits(stealNet_io_connSS_0_data_availableTask_bits),
    .io_connSS_0_data_qOutTask_ready(stealNet_io_connSS_0_data_qOutTask_ready),
    .io_connSS_0_data_qOutTask_valid(stealNet_io_connSS_0_data_qOutTask_valid),
    .io_connSS_0_data_qOutTask_bits(stealNet_io_connSS_0_data_qOutTask_bits),
    .io_connSS_1_ctrl_serveStealReq_ready(stealNet_io_connSS_1_ctrl_serveStealReq_ready),
    .io_connSS_1_ctrl_serveStealReq_valid(stealNet_io_connSS_1_ctrl_serveStealReq_valid),
    .io_connSS_1_data_qOutTask_ready(stealNet_io_connSS_1_data_qOutTask_ready),
    .io_connSS_1_data_qOutTask_valid(stealNet_io_connSS_1_data_qOutTask_valid),
    .io_connSS_1_data_qOutTask_bits(stealNet_io_connSS_1_data_qOutTask_bits),
    .io_connSS_2_ctrl_serveStealReq_ready(stealNet_io_connSS_2_ctrl_serveStealReq_ready),
    .io_connSS_2_ctrl_serveStealReq_valid(stealNet_io_connSS_2_ctrl_serveStealReq_valid),
    .io_connSS_2_data_qOutTask_ready(stealNet_io_connSS_2_data_qOutTask_ready),
    .io_connSS_2_data_qOutTask_valid(stealNet_io_connSS_2_data_qOutTask_valid),
    .io_connSS_2_data_qOutTask_bits(stealNet_io_connSS_2_data_qOutTask_bits),
    .io_connSS_3_ctrl_serveStealReq_ready(stealNet_io_connSS_3_ctrl_serveStealReq_ready),
    .io_connSS_3_ctrl_serveStealReq_valid(stealNet_io_connSS_3_ctrl_serveStealReq_valid),
    .io_connSS_3_ctrl_stealReq_ready(stealNet_io_connSS_3_ctrl_stealReq_ready),
    .io_connSS_3_ctrl_stealReq_valid(stealNet_io_connSS_3_ctrl_stealReq_valid),
    .io_connSS_3_data_availableTask_ready(stealNet_io_connSS_3_data_availableTask_ready),
    .io_connSS_3_data_availableTask_valid(stealNet_io_connSS_3_data_availableTask_valid),
    .io_connSS_3_data_availableTask_bits(stealNet_io_connSS_3_data_availableTask_bits),
    .io_connSS_3_data_qOutTask_ready(stealNet_io_connSS_3_data_qOutTask_ready),
    .io_connSS_3_data_qOutTask_valid(stealNet_io_connSS_3_data_qOutTask_valid),
    .io_connSS_3_data_qOutTask_bits(stealNet_io_connSS_3_data_qOutTask_bits),
    .io_connSS_4_ctrl_serveStealReq_ready(stealNet_io_connSS_4_ctrl_serveStealReq_ready),
    .io_connSS_4_ctrl_serveStealReq_valid(stealNet_io_connSS_4_ctrl_serveStealReq_valid),
    .io_connSS_4_ctrl_stealReq_ready(stealNet_io_connSS_4_ctrl_stealReq_ready),
    .io_connSS_4_ctrl_stealReq_valid(stealNet_io_connSS_4_ctrl_stealReq_valid),
    .io_connSS_4_data_availableTask_ready(stealNet_io_connSS_4_data_availableTask_ready),
    .io_connSS_4_data_availableTask_valid(stealNet_io_connSS_4_data_availableTask_valid),
    .io_connSS_4_data_availableTask_bits(stealNet_io_connSS_4_data_availableTask_bits),
    .io_connSS_4_data_qOutTask_ready(stealNet_io_connSS_4_data_qOutTask_ready),
    .io_connSS_4_data_qOutTask_valid(stealNet_io_connSS_4_data_qOutTask_valid),
    .io_connSS_4_data_qOutTask_bits(stealNet_io_connSS_4_data_qOutTask_bits),
    .io_connSS_5_ctrl_serveStealReq_ready(stealNet_io_connSS_5_ctrl_serveStealReq_ready),
    .io_connSS_5_ctrl_serveStealReq_valid(stealNet_io_connSS_5_ctrl_serveStealReq_valid),
    .io_connSS_5_ctrl_stealReq_ready(stealNet_io_connSS_5_ctrl_stealReq_ready),
    .io_connSS_5_ctrl_stealReq_valid(stealNet_io_connSS_5_ctrl_stealReq_valid),
    .io_connSS_5_data_availableTask_ready(stealNet_io_connSS_5_data_availableTask_ready),
    .io_connSS_5_data_availableTask_valid(stealNet_io_connSS_5_data_availableTask_valid),
    .io_connSS_5_data_availableTask_bits(stealNet_io_connSS_5_data_availableTask_bits),
    .io_connSS_5_data_qOutTask_ready(stealNet_io_connSS_5_data_qOutTask_ready),
    .io_connSS_5_data_qOutTask_valid(stealNet_io_connSS_5_data_qOutTask_valid),
    .io_connSS_5_data_qOutTask_bits(stealNet_io_connSS_5_data_qOutTask_bits),
    .io_connSS_6_ctrl_serveStealReq_ready(stealNet_io_connSS_6_ctrl_serveStealReq_ready),
    .io_connSS_6_ctrl_serveStealReq_valid(stealNet_io_connSS_6_ctrl_serveStealReq_valid),
    .io_connSS_6_ctrl_stealReq_ready(stealNet_io_connSS_6_ctrl_stealReq_ready),
    .io_connSS_6_ctrl_stealReq_valid(stealNet_io_connSS_6_ctrl_stealReq_valid),
    .io_connSS_6_data_availableTask_ready(stealNet_io_connSS_6_data_availableTask_ready),
    .io_connSS_6_data_availableTask_valid(stealNet_io_connSS_6_data_availableTask_valid),
    .io_connSS_6_data_availableTask_bits(stealNet_io_connSS_6_data_availableTask_bits),
    .io_connSS_6_data_qOutTask_ready(stealNet_io_connSS_6_data_qOutTask_ready),
    .io_connSS_6_data_qOutTask_valid(stealNet_io_connSS_6_data_qOutTask_valid),
    .io_connSS_6_data_qOutTask_bits(stealNet_io_connSS_6_data_qOutTask_bits),
    .io_connSS_7_ctrl_serveStealReq_ready(stealNet_io_connSS_7_ctrl_serveStealReq_ready),
    .io_connSS_7_ctrl_serveStealReq_valid(stealNet_io_connSS_7_ctrl_serveStealReq_valid),
    .io_connSS_7_ctrl_stealReq_ready(stealNet_io_connSS_7_ctrl_stealReq_ready),
    .io_connSS_7_ctrl_stealReq_valid(stealNet_io_connSS_7_ctrl_stealReq_valid),
    .io_connSS_7_data_availableTask_ready(stealNet_io_connSS_7_data_availableTask_ready),
    .io_connSS_7_data_availableTask_valid(stealNet_io_connSS_7_data_availableTask_valid),
    .io_connSS_7_data_availableTask_bits(stealNet_io_connSS_7_data_availableTask_bits),
    .io_connSS_7_data_qOutTask_ready(stealNet_io_connSS_7_data_qOutTask_ready),
    .io_connSS_7_data_qOutTask_valid(stealNet_io_connSS_7_data_qOutTask_valid),
    .io_connSS_7_data_qOutTask_bits(stealNet_io_connSS_7_data_qOutTask_bits),
    .io_connSS_8_ctrl_serveStealReq_ready(stealNet_io_connSS_8_ctrl_serveStealReq_ready),
    .io_connSS_8_ctrl_serveStealReq_valid(stealNet_io_connSS_8_ctrl_serveStealReq_valid),
    .io_connSS_8_ctrl_stealReq_ready(stealNet_io_connSS_8_ctrl_stealReq_ready),
    .io_connSS_8_ctrl_stealReq_valid(stealNet_io_connSS_8_ctrl_stealReq_valid),
    .io_connSS_8_data_availableTask_ready(stealNet_io_connSS_8_data_availableTask_ready),
    .io_connSS_8_data_availableTask_valid(stealNet_io_connSS_8_data_availableTask_valid),
    .io_connSS_8_data_availableTask_bits(stealNet_io_connSS_8_data_availableTask_bits),
    .io_connSS_8_data_qOutTask_ready(stealNet_io_connSS_8_data_qOutTask_ready),
    .io_connSS_8_data_qOutTask_valid(stealNet_io_connSS_8_data_qOutTask_valid),
    .io_connSS_8_data_qOutTask_bits(stealNet_io_connSS_8_data_qOutTask_bits),
    .io_connSS_9_ctrl_serveStealReq_ready(stealNet_io_connSS_9_ctrl_serveStealReq_ready),
    .io_connSS_9_ctrl_serveStealReq_valid(stealNet_io_connSS_9_ctrl_serveStealReq_valid),
    .io_connSS_9_ctrl_stealReq_ready(stealNet_io_connSS_9_ctrl_stealReq_ready),
    .io_connSS_9_ctrl_stealReq_valid(stealNet_io_connSS_9_ctrl_stealReq_valid),
    .io_connSS_9_data_availableTask_ready(stealNet_io_connSS_9_data_availableTask_ready),
    .io_connSS_9_data_availableTask_valid(stealNet_io_connSS_9_data_availableTask_valid),
    .io_connSS_9_data_availableTask_bits(stealNet_io_connSS_9_data_availableTask_bits),
    .io_connSS_9_data_qOutTask_ready(stealNet_io_connSS_9_data_qOutTask_ready),
    .io_connSS_9_data_qOutTask_valid(stealNet_io_connSS_9_data_qOutTask_valid),
    .io_connSS_9_data_qOutTask_bits(stealNet_io_connSS_9_data_qOutTask_bits),
    .io_connSS_10_ctrl_serveStealReq_ready(stealNet_io_connSS_10_ctrl_serveStealReq_ready),
    .io_connSS_10_ctrl_serveStealReq_valid(stealNet_io_connSS_10_ctrl_serveStealReq_valid),
    .io_connSS_10_ctrl_stealReq_ready(stealNet_io_connSS_10_ctrl_stealReq_ready),
    .io_connSS_10_ctrl_stealReq_valid(stealNet_io_connSS_10_ctrl_stealReq_valid),
    .io_connSS_10_data_availableTask_ready(stealNet_io_connSS_10_data_availableTask_ready),
    .io_connSS_10_data_availableTask_valid(stealNet_io_connSS_10_data_availableTask_valid),
    .io_connSS_10_data_availableTask_bits(stealNet_io_connSS_10_data_availableTask_bits),
    .io_connSS_10_data_qOutTask_ready(stealNet_io_connSS_10_data_qOutTask_ready),
    .io_connSS_10_data_qOutTask_valid(stealNet_io_connSS_10_data_qOutTask_valid),
    .io_connSS_10_data_qOutTask_bits(stealNet_io_connSS_10_data_qOutTask_bits),
    .io_connSS_11_ctrl_serveStealReq_ready(stealNet_io_connSS_11_ctrl_serveStealReq_ready),
    .io_connSS_11_ctrl_serveStealReq_valid(stealNet_io_connSS_11_ctrl_serveStealReq_valid),
    .io_connSS_11_ctrl_stealReq_ready(stealNet_io_connSS_11_ctrl_stealReq_ready),
    .io_connSS_11_ctrl_stealReq_valid(stealNet_io_connSS_11_ctrl_stealReq_valid),
    .io_connSS_11_data_availableTask_ready(stealNet_io_connSS_11_data_availableTask_ready),
    .io_connSS_11_data_availableTask_valid(stealNet_io_connSS_11_data_availableTask_valid),
    .io_connSS_11_data_availableTask_bits(stealNet_io_connSS_11_data_availableTask_bits),
    .io_connSS_11_data_qOutTask_ready(stealNet_io_connSS_11_data_qOutTask_ready),
    .io_connSS_11_data_qOutTask_valid(stealNet_io_connSS_11_data_qOutTask_valid),
    .io_connSS_11_data_qOutTask_bits(stealNet_io_connSS_11_data_qOutTask_bits),
    .io_connSS_12_ctrl_serveStealReq_ready(stealNet_io_connSS_12_ctrl_serveStealReq_ready),
    .io_connSS_12_ctrl_serveStealReq_valid(stealNet_io_connSS_12_ctrl_serveStealReq_valid),
    .io_connSS_12_ctrl_stealReq_ready(stealNet_io_connSS_12_ctrl_stealReq_ready),
    .io_connSS_12_ctrl_stealReq_valid(stealNet_io_connSS_12_ctrl_stealReq_valid),
    .io_connSS_12_data_availableTask_ready(stealNet_io_connSS_12_data_availableTask_ready),
    .io_connSS_12_data_availableTask_valid(stealNet_io_connSS_12_data_availableTask_valid),
    .io_connSS_12_data_availableTask_bits(stealNet_io_connSS_12_data_availableTask_bits),
    .io_connSS_12_data_qOutTask_ready(stealNet_io_connSS_12_data_qOutTask_ready),
    .io_connSS_12_data_qOutTask_valid(stealNet_io_connSS_12_data_qOutTask_valid),
    .io_connSS_12_data_qOutTask_bits(stealNet_io_connSS_12_data_qOutTask_bits),
    .io_connSS_13_ctrl_serveStealReq_ready(stealNet_io_connSS_13_ctrl_serveStealReq_ready),
    .io_connSS_13_ctrl_serveStealReq_valid(stealNet_io_connSS_13_ctrl_serveStealReq_valid),
    .io_connSS_13_ctrl_stealReq_ready(stealNet_io_connSS_13_ctrl_stealReq_ready),
    .io_connSS_13_ctrl_stealReq_valid(stealNet_io_connSS_13_ctrl_stealReq_valid),
    .io_connSS_13_data_availableTask_ready(stealNet_io_connSS_13_data_availableTask_ready),
    .io_connSS_13_data_availableTask_valid(stealNet_io_connSS_13_data_availableTask_valid),
    .io_connSS_13_data_availableTask_bits(stealNet_io_connSS_13_data_availableTask_bits),
    .io_connSS_13_data_qOutTask_ready(stealNet_io_connSS_13_data_qOutTask_ready),
    .io_connSS_13_data_qOutTask_valid(stealNet_io_connSS_13_data_qOutTask_valid),
    .io_connSS_13_data_qOutTask_bits(stealNet_io_connSS_13_data_qOutTask_bits),
    .io_connSS_14_ctrl_serveStealReq_ready(stealNet_io_connSS_14_ctrl_serveStealReq_ready),
    .io_connSS_14_ctrl_serveStealReq_valid(stealNet_io_connSS_14_ctrl_serveStealReq_valid),
    .io_connSS_14_ctrl_stealReq_ready(stealNet_io_connSS_14_ctrl_stealReq_ready),
    .io_connSS_14_ctrl_stealReq_valid(stealNet_io_connSS_14_ctrl_stealReq_valid),
    .io_connSS_14_data_availableTask_ready(stealNet_io_connSS_14_data_availableTask_ready),
    .io_connSS_14_data_availableTask_valid(stealNet_io_connSS_14_data_availableTask_valid),
    .io_connSS_14_data_availableTask_bits(stealNet_io_connSS_14_data_availableTask_bits),
    .io_connSS_14_data_qOutTask_ready(stealNet_io_connSS_14_data_qOutTask_ready),
    .io_connSS_14_data_qOutTask_valid(stealNet_io_connSS_14_data_qOutTask_valid),
    .io_connSS_14_data_qOutTask_bits(stealNet_io_connSS_14_data_qOutTask_bits),
    .io_connSS_15_ctrl_serveStealReq_ready(stealNet_io_connSS_15_ctrl_serveStealReq_ready),
    .io_connSS_15_ctrl_serveStealReq_valid(stealNet_io_connSS_15_ctrl_serveStealReq_valid),
    .io_connSS_15_ctrl_stealReq_ready(stealNet_io_connSS_15_ctrl_stealReq_ready),
    .io_connSS_15_ctrl_stealReq_valid(stealNet_io_connSS_15_ctrl_stealReq_valid),
    .io_connSS_15_data_availableTask_ready(stealNet_io_connSS_15_data_availableTask_ready),
    .io_connSS_15_data_availableTask_valid(stealNet_io_connSS_15_data_availableTask_valid),
    .io_connSS_15_data_availableTask_bits(stealNet_io_connSS_15_data_availableTask_bits),
    .io_connSS_15_data_qOutTask_ready(stealNet_io_connSS_15_data_qOutTask_ready),
    .io_connSS_15_data_qOutTask_valid(stealNet_io_connSS_15_data_qOutTask_valid),
    .io_connSS_15_data_qOutTask_bits(stealNet_io_connSS_15_data_qOutTask_bits),
    .io_connSS_16_ctrl_serveStealReq_ready(stealNet_io_connSS_16_ctrl_serveStealReq_ready),
    .io_connSS_16_ctrl_serveStealReq_valid(stealNet_io_connSS_16_ctrl_serveStealReq_valid),
    .io_connSS_16_ctrl_stealReq_ready(stealNet_io_connSS_16_ctrl_stealReq_ready),
    .io_connSS_16_ctrl_stealReq_valid(stealNet_io_connSS_16_ctrl_stealReq_valid),
    .io_connSS_16_data_availableTask_ready(stealNet_io_connSS_16_data_availableTask_ready),
    .io_connSS_16_data_availableTask_valid(stealNet_io_connSS_16_data_availableTask_valid),
    .io_connSS_16_data_availableTask_bits(stealNet_io_connSS_16_data_availableTask_bits),
    .io_connSS_16_data_qOutTask_ready(stealNet_io_connSS_16_data_qOutTask_ready),
    .io_connSS_16_data_qOutTask_valid(stealNet_io_connSS_16_data_qOutTask_valid),
    .io_connSS_16_data_qOutTask_bits(stealNet_io_connSS_16_data_qOutTask_bits),
    .io_connSS_17_ctrl_serveStealReq_ready(stealNet_io_connSS_17_ctrl_serveStealReq_ready),
    .io_connSS_17_ctrl_serveStealReq_valid(stealNet_io_connSS_17_ctrl_serveStealReq_valid),
    .io_connSS_17_ctrl_stealReq_ready(stealNet_io_connSS_17_ctrl_stealReq_ready),
    .io_connSS_17_ctrl_stealReq_valid(stealNet_io_connSS_17_ctrl_stealReq_valid),
    .io_connSS_17_data_availableTask_ready(stealNet_io_connSS_17_data_availableTask_ready),
    .io_connSS_17_data_availableTask_valid(stealNet_io_connSS_17_data_availableTask_valid),
    .io_connSS_17_data_availableTask_bits(stealNet_io_connSS_17_data_availableTask_bits),
    .io_connSS_17_data_qOutTask_ready(stealNet_io_connSS_17_data_qOutTask_ready),
    .io_connSS_17_data_qOutTask_valid(stealNet_io_connSS_17_data_qOutTask_valid),
    .io_connSS_17_data_qOutTask_bits(stealNet_io_connSS_17_data_qOutTask_bits),
    .io_connSS_18_ctrl_serveStealReq_ready(stealNet_io_connSS_18_ctrl_serveStealReq_ready),
    .io_connSS_18_ctrl_serveStealReq_valid(stealNet_io_connSS_18_ctrl_serveStealReq_valid),
    .io_connSS_18_ctrl_stealReq_ready(stealNet_io_connSS_18_ctrl_stealReq_ready),
    .io_connSS_18_ctrl_stealReq_valid(stealNet_io_connSS_18_ctrl_stealReq_valid),
    .io_connSS_18_data_availableTask_ready(stealNet_io_connSS_18_data_availableTask_ready),
    .io_connSS_18_data_availableTask_valid(stealNet_io_connSS_18_data_availableTask_valid),
    .io_connSS_18_data_availableTask_bits(stealNet_io_connSS_18_data_availableTask_bits),
    .io_connSS_18_data_qOutTask_ready(stealNet_io_connSS_18_data_qOutTask_ready),
    .io_connSS_18_data_qOutTask_valid(stealNet_io_connSS_18_data_qOutTask_valid),
    .io_connSS_18_data_qOutTask_bits(stealNet_io_connSS_18_data_qOutTask_bits),
    .io_connSS_19_ctrl_serveStealReq_ready(stealNet_io_connSS_19_ctrl_serveStealReq_ready),
    .io_connSS_19_ctrl_serveStealReq_valid(stealNet_io_connSS_19_ctrl_serveStealReq_valid),
    .io_connSS_19_ctrl_stealReq_ready(stealNet_io_connSS_19_ctrl_stealReq_ready),
    .io_connSS_19_ctrl_stealReq_valid(stealNet_io_connSS_19_ctrl_stealReq_valid),
    .io_connSS_19_data_availableTask_ready(stealNet_io_connSS_19_data_availableTask_ready),
    .io_connSS_19_data_availableTask_valid(stealNet_io_connSS_19_data_availableTask_valid),
    .io_connSS_19_data_availableTask_bits(stealNet_io_connSS_19_data_availableTask_bits),
    .io_connSS_19_data_qOutTask_ready(stealNet_io_connSS_19_data_qOutTask_ready),
    .io_connSS_19_data_qOutTask_valid(stealNet_io_connSS_19_data_qOutTask_valid),
    .io_connSS_19_data_qOutTask_bits(stealNet_io_connSS_19_data_qOutTask_bits),
    .io_connSS_20_ctrl_serveStealReq_ready(stealNet_io_connSS_20_ctrl_serveStealReq_ready),
    .io_connSS_20_ctrl_serveStealReq_valid(stealNet_io_connSS_20_ctrl_serveStealReq_valid),
    .io_connSS_20_ctrl_stealReq_ready(stealNet_io_connSS_20_ctrl_stealReq_ready),
    .io_connSS_20_ctrl_stealReq_valid(stealNet_io_connSS_20_ctrl_stealReq_valid),
    .io_connSS_20_data_availableTask_ready(stealNet_io_connSS_20_data_availableTask_ready),
    .io_connSS_20_data_availableTask_valid(stealNet_io_connSS_20_data_availableTask_valid),
    .io_connSS_20_data_availableTask_bits(stealNet_io_connSS_20_data_availableTask_bits),
    .io_connSS_20_data_qOutTask_ready(stealNet_io_connSS_20_data_qOutTask_ready),
    .io_connSS_20_data_qOutTask_valid(stealNet_io_connSS_20_data_qOutTask_valid),
    .io_connSS_20_data_qOutTask_bits(stealNet_io_connSS_20_data_qOutTask_bits),
    .io_connSS_21_ctrl_serveStealReq_ready(stealNet_io_connSS_21_ctrl_serveStealReq_ready),
    .io_connSS_21_ctrl_serveStealReq_valid(stealNet_io_connSS_21_ctrl_serveStealReq_valid),
    .io_connSS_21_ctrl_stealReq_ready(stealNet_io_connSS_21_ctrl_stealReq_ready),
    .io_connSS_21_ctrl_stealReq_valid(stealNet_io_connSS_21_ctrl_stealReq_valid),
    .io_connSS_21_data_availableTask_ready(stealNet_io_connSS_21_data_availableTask_ready),
    .io_connSS_21_data_availableTask_valid(stealNet_io_connSS_21_data_availableTask_valid),
    .io_connSS_21_data_availableTask_bits(stealNet_io_connSS_21_data_availableTask_bits),
    .io_connSS_21_data_qOutTask_ready(stealNet_io_connSS_21_data_qOutTask_ready),
    .io_connSS_21_data_qOutTask_valid(stealNet_io_connSS_21_data_qOutTask_valid),
    .io_connSS_21_data_qOutTask_bits(stealNet_io_connSS_21_data_qOutTask_bits),
    .io_connSS_22_ctrl_serveStealReq_ready(stealNet_io_connSS_22_ctrl_serveStealReq_ready),
    .io_connSS_22_ctrl_serveStealReq_valid(stealNet_io_connSS_22_ctrl_serveStealReq_valid),
    .io_connSS_22_ctrl_stealReq_ready(stealNet_io_connSS_22_ctrl_stealReq_ready),
    .io_connSS_22_ctrl_stealReq_valid(stealNet_io_connSS_22_ctrl_stealReq_valid),
    .io_connSS_22_data_availableTask_ready(stealNet_io_connSS_22_data_availableTask_ready),
    .io_connSS_22_data_availableTask_valid(stealNet_io_connSS_22_data_availableTask_valid),
    .io_connSS_22_data_availableTask_bits(stealNet_io_connSS_22_data_availableTask_bits),
    .io_connSS_22_data_qOutTask_ready(stealNet_io_connSS_22_data_qOutTask_ready),
    .io_connSS_22_data_qOutTask_valid(stealNet_io_connSS_22_data_qOutTask_valid),
    .io_connSS_22_data_qOutTask_bits(stealNet_io_connSS_22_data_qOutTask_bits),
    .io_connSS_23_ctrl_serveStealReq_ready(stealNet_io_connSS_23_ctrl_serveStealReq_ready),
    .io_connSS_23_ctrl_serveStealReq_valid(stealNet_io_connSS_23_ctrl_serveStealReq_valid),
    .io_connSS_23_ctrl_stealReq_ready(stealNet_io_connSS_23_ctrl_stealReq_ready),
    .io_connSS_23_ctrl_stealReq_valid(stealNet_io_connSS_23_ctrl_stealReq_valid),
    .io_connSS_23_data_availableTask_ready(stealNet_io_connSS_23_data_availableTask_ready),
    .io_connSS_23_data_availableTask_valid(stealNet_io_connSS_23_data_availableTask_valid),
    .io_connSS_23_data_availableTask_bits(stealNet_io_connSS_23_data_availableTask_bits),
    .io_connSS_23_data_qOutTask_ready(stealNet_io_connSS_23_data_qOutTask_ready),
    .io_connSS_23_data_qOutTask_valid(stealNet_io_connSS_23_data_qOutTask_valid),
    .io_connSS_23_data_qOutTask_bits(stealNet_io_connSS_23_data_qOutTask_bits),
    .io_connSS_24_ctrl_serveStealReq_ready(stealNet_io_connSS_24_ctrl_serveStealReq_ready),
    .io_connSS_24_ctrl_serveStealReq_valid(stealNet_io_connSS_24_ctrl_serveStealReq_valid),
    .io_connSS_24_ctrl_stealReq_ready(stealNet_io_connSS_24_ctrl_stealReq_ready),
    .io_connSS_24_ctrl_stealReq_valid(stealNet_io_connSS_24_ctrl_stealReq_valid),
    .io_connSS_24_data_availableTask_ready(stealNet_io_connSS_24_data_availableTask_ready),
    .io_connSS_24_data_availableTask_valid(stealNet_io_connSS_24_data_availableTask_valid),
    .io_connSS_24_data_availableTask_bits(stealNet_io_connSS_24_data_availableTask_bits),
    .io_connSS_24_data_qOutTask_ready(stealNet_io_connSS_24_data_qOutTask_ready),
    .io_connSS_24_data_qOutTask_valid(stealNet_io_connSS_24_data_qOutTask_valid),
    .io_connSS_24_data_qOutTask_bits(stealNet_io_connSS_24_data_qOutTask_bits),
    .io_connSS_25_ctrl_serveStealReq_ready(stealNet_io_connSS_25_ctrl_serveStealReq_ready),
    .io_connSS_25_ctrl_serveStealReq_valid(stealNet_io_connSS_25_ctrl_serveStealReq_valid),
    .io_connSS_25_ctrl_stealReq_ready(stealNet_io_connSS_25_ctrl_stealReq_ready),
    .io_connSS_25_ctrl_stealReq_valid(stealNet_io_connSS_25_ctrl_stealReq_valid),
    .io_connSS_25_data_availableTask_ready(stealNet_io_connSS_25_data_availableTask_ready),
    .io_connSS_25_data_availableTask_valid(stealNet_io_connSS_25_data_availableTask_valid),
    .io_connSS_25_data_availableTask_bits(stealNet_io_connSS_25_data_availableTask_bits),
    .io_connSS_25_data_qOutTask_ready(stealNet_io_connSS_25_data_qOutTask_ready),
    .io_connSS_25_data_qOutTask_valid(stealNet_io_connSS_25_data_qOutTask_valid),
    .io_connSS_25_data_qOutTask_bits(stealNet_io_connSS_25_data_qOutTask_bits),
    .io_connSS_26_ctrl_serveStealReq_ready(stealNet_io_connSS_26_ctrl_serveStealReq_ready),
    .io_connSS_26_ctrl_serveStealReq_valid(stealNet_io_connSS_26_ctrl_serveStealReq_valid),
    .io_connSS_26_ctrl_stealReq_ready(stealNet_io_connSS_26_ctrl_stealReq_ready),
    .io_connSS_26_ctrl_stealReq_valid(stealNet_io_connSS_26_ctrl_stealReq_valid),
    .io_connSS_26_data_availableTask_ready(stealNet_io_connSS_26_data_availableTask_ready),
    .io_connSS_26_data_availableTask_valid(stealNet_io_connSS_26_data_availableTask_valid),
    .io_connSS_26_data_availableTask_bits(stealNet_io_connSS_26_data_availableTask_bits),
    .io_connSS_26_data_qOutTask_ready(stealNet_io_connSS_26_data_qOutTask_ready),
    .io_connSS_26_data_qOutTask_valid(stealNet_io_connSS_26_data_qOutTask_valid),
    .io_connSS_26_data_qOutTask_bits(stealNet_io_connSS_26_data_qOutTask_bits),
    .io_connSS_27_ctrl_serveStealReq_ready(stealNet_io_connSS_27_ctrl_serveStealReq_ready),
    .io_connSS_27_ctrl_serveStealReq_valid(stealNet_io_connSS_27_ctrl_serveStealReq_valid),
    .io_connSS_27_ctrl_stealReq_ready(stealNet_io_connSS_27_ctrl_stealReq_ready),
    .io_connSS_27_ctrl_stealReq_valid(stealNet_io_connSS_27_ctrl_stealReq_valid),
    .io_connSS_27_data_availableTask_ready(stealNet_io_connSS_27_data_availableTask_ready),
    .io_connSS_27_data_availableTask_valid(stealNet_io_connSS_27_data_availableTask_valid),
    .io_connSS_27_data_availableTask_bits(stealNet_io_connSS_27_data_availableTask_bits),
    .io_connSS_27_data_qOutTask_ready(stealNet_io_connSS_27_data_qOutTask_ready),
    .io_connSS_27_data_qOutTask_valid(stealNet_io_connSS_27_data_qOutTask_valid),
    .io_connSS_27_data_qOutTask_bits(stealNet_io_connSS_27_data_qOutTask_bits),
    .io_connSS_28_ctrl_serveStealReq_ready(stealNet_io_connSS_28_ctrl_serveStealReq_ready),
    .io_connSS_28_ctrl_serveStealReq_valid(stealNet_io_connSS_28_ctrl_serveStealReq_valid),
    .io_connSS_28_ctrl_stealReq_ready(stealNet_io_connSS_28_ctrl_stealReq_ready),
    .io_connSS_28_ctrl_stealReq_valid(stealNet_io_connSS_28_ctrl_stealReq_valid),
    .io_connSS_28_data_availableTask_ready(stealNet_io_connSS_28_data_availableTask_ready),
    .io_connSS_28_data_availableTask_valid(stealNet_io_connSS_28_data_availableTask_valid),
    .io_connSS_28_data_availableTask_bits(stealNet_io_connSS_28_data_availableTask_bits),
    .io_connSS_28_data_qOutTask_ready(stealNet_io_connSS_28_data_qOutTask_ready),
    .io_connSS_28_data_qOutTask_valid(stealNet_io_connSS_28_data_qOutTask_valid),
    .io_connSS_28_data_qOutTask_bits(stealNet_io_connSS_28_data_qOutTask_bits),
    .io_connSS_29_ctrl_serveStealReq_ready(stealNet_io_connSS_29_ctrl_serveStealReq_ready),
    .io_connSS_29_ctrl_serveStealReq_valid(stealNet_io_connSS_29_ctrl_serveStealReq_valid),
    .io_connSS_29_ctrl_stealReq_ready(stealNet_io_connSS_29_ctrl_stealReq_ready),
    .io_connSS_29_ctrl_stealReq_valid(stealNet_io_connSS_29_ctrl_stealReq_valid),
    .io_connSS_29_data_availableTask_ready(stealNet_io_connSS_29_data_availableTask_ready),
    .io_connSS_29_data_availableTask_valid(stealNet_io_connSS_29_data_availableTask_valid),
    .io_connSS_29_data_availableTask_bits(stealNet_io_connSS_29_data_availableTask_bits),
    .io_connSS_29_data_qOutTask_ready(stealNet_io_connSS_29_data_qOutTask_ready),
    .io_connSS_29_data_qOutTask_valid(stealNet_io_connSS_29_data_qOutTask_valid),
    .io_connSS_29_data_qOutTask_bits(stealNet_io_connSS_29_data_qOutTask_bits),
    .io_connSS_30_ctrl_serveStealReq_ready(stealNet_io_connSS_30_ctrl_serveStealReq_ready),
    .io_connSS_30_ctrl_serveStealReq_valid(stealNet_io_connSS_30_ctrl_serveStealReq_valid),
    .io_connSS_30_ctrl_stealReq_ready(stealNet_io_connSS_30_ctrl_stealReq_ready),
    .io_connSS_30_ctrl_stealReq_valid(stealNet_io_connSS_30_ctrl_stealReq_valid),
    .io_connSS_30_data_availableTask_ready(stealNet_io_connSS_30_data_availableTask_ready),
    .io_connSS_30_data_availableTask_valid(stealNet_io_connSS_30_data_availableTask_valid),
    .io_connSS_30_data_availableTask_bits(stealNet_io_connSS_30_data_availableTask_bits),
    .io_connSS_30_data_qOutTask_ready(stealNet_io_connSS_30_data_qOutTask_ready),
    .io_connSS_30_data_qOutTask_valid(stealNet_io_connSS_30_data_qOutTask_valid),
    .io_connSS_30_data_qOutTask_bits(stealNet_io_connSS_30_data_qOutTask_bits),
    .io_connSS_31_ctrl_serveStealReq_ready(stealNet_io_connSS_31_ctrl_serveStealReq_ready),
    .io_connSS_31_ctrl_serveStealReq_valid(stealNet_io_connSS_31_ctrl_serveStealReq_valid),
    .io_connSS_31_ctrl_stealReq_ready(stealNet_io_connSS_31_ctrl_stealReq_ready),
    .io_connSS_31_ctrl_stealReq_valid(stealNet_io_connSS_31_ctrl_stealReq_valid),
    .io_connSS_31_data_availableTask_ready(stealNet_io_connSS_31_data_availableTask_ready),
    .io_connSS_31_data_availableTask_valid(stealNet_io_connSS_31_data_availableTask_valid),
    .io_connSS_31_data_availableTask_bits(stealNet_io_connSS_31_data_availableTask_bits),
    .io_connSS_31_data_qOutTask_ready(stealNet_io_connSS_31_data_qOutTask_ready),
    .io_connSS_31_data_qOutTask_valid(stealNet_io_connSS_31_data_qOutTask_valid),
    .io_connSS_31_data_qOutTask_bits(stealNet_io_connSS_31_data_qOutTask_bits),
    .io_connSS_32_ctrl_serveStealReq_ready(stealNet_io_connSS_32_ctrl_serveStealReq_ready),
    .io_connSS_32_ctrl_serveStealReq_valid(stealNet_io_connSS_32_ctrl_serveStealReq_valid),
    .io_connSS_32_ctrl_stealReq_ready(stealNet_io_connSS_32_ctrl_stealReq_ready),
    .io_connSS_32_ctrl_stealReq_valid(stealNet_io_connSS_32_ctrl_stealReq_valid),
    .io_connSS_32_data_availableTask_ready(stealNet_io_connSS_32_data_availableTask_ready),
    .io_connSS_32_data_availableTask_valid(stealNet_io_connSS_32_data_availableTask_valid),
    .io_connSS_32_data_availableTask_bits(stealNet_io_connSS_32_data_availableTask_bits),
    .io_connSS_32_data_qOutTask_ready(stealNet_io_connSS_32_data_qOutTask_ready),
    .io_connSS_32_data_qOutTask_valid(stealNet_io_connSS_32_data_qOutTask_valid),
    .io_connSS_32_data_qOutTask_bits(stealNet_io_connSS_32_data_qOutTask_bits),
    .io_connSS_33_ctrl_serveStealReq_ready(stealNet_io_connSS_33_ctrl_serveStealReq_ready),
    .io_connSS_33_ctrl_serveStealReq_valid(stealNet_io_connSS_33_ctrl_serveStealReq_valid),
    .io_connSS_33_ctrl_stealReq_ready(stealNet_io_connSS_33_ctrl_stealReq_ready),
    .io_connSS_33_ctrl_stealReq_valid(stealNet_io_connSS_33_ctrl_stealReq_valid),
    .io_connSS_33_data_availableTask_ready(stealNet_io_connSS_33_data_availableTask_ready),
    .io_connSS_33_data_availableTask_valid(stealNet_io_connSS_33_data_availableTask_valid),
    .io_connSS_33_data_availableTask_bits(stealNet_io_connSS_33_data_availableTask_bits),
    .io_connSS_33_data_qOutTask_ready(stealNet_io_connSS_33_data_qOutTask_ready),
    .io_connSS_33_data_qOutTask_valid(stealNet_io_connSS_33_data_qOutTask_valid),
    .io_connSS_33_data_qOutTask_bits(stealNet_io_connSS_33_data_qOutTask_bits),
    .io_connSS_34_ctrl_serveStealReq_ready(stealNet_io_connSS_34_ctrl_serveStealReq_ready),
    .io_connSS_34_ctrl_serveStealReq_valid(stealNet_io_connSS_34_ctrl_serveStealReq_valid),
    .io_connSS_34_ctrl_stealReq_ready(stealNet_io_connSS_34_ctrl_stealReq_ready),
    .io_connSS_34_ctrl_stealReq_valid(stealNet_io_connSS_34_ctrl_stealReq_valid),
    .io_connSS_34_data_availableTask_ready(stealNet_io_connSS_34_data_availableTask_ready),
    .io_connSS_34_data_availableTask_valid(stealNet_io_connSS_34_data_availableTask_valid),
    .io_connSS_34_data_availableTask_bits(stealNet_io_connSS_34_data_availableTask_bits),
    .io_connSS_34_data_qOutTask_ready(stealNet_io_connSS_34_data_qOutTask_ready),
    .io_connSS_34_data_qOutTask_valid(stealNet_io_connSS_34_data_qOutTask_valid),
    .io_connSS_34_data_qOutTask_bits(stealNet_io_connSS_34_data_qOutTask_bits),
    .io_connSS_35_ctrl_serveStealReq_ready(stealNet_io_connSS_35_ctrl_serveStealReq_ready),
    .io_connSS_35_ctrl_serveStealReq_valid(stealNet_io_connSS_35_ctrl_serveStealReq_valid),
    .io_connSS_35_ctrl_stealReq_ready(stealNet_io_connSS_35_ctrl_stealReq_ready),
    .io_connSS_35_ctrl_stealReq_valid(stealNet_io_connSS_35_ctrl_stealReq_valid),
    .io_connSS_35_data_availableTask_ready(stealNet_io_connSS_35_data_availableTask_ready),
    .io_connSS_35_data_availableTask_valid(stealNet_io_connSS_35_data_availableTask_valid),
    .io_connSS_35_data_availableTask_bits(stealNet_io_connSS_35_data_availableTask_bits),
    .io_connSS_35_data_qOutTask_ready(stealNet_io_connSS_35_data_qOutTask_ready),
    .io_connSS_35_data_qOutTask_valid(stealNet_io_connSS_35_data_qOutTask_valid),
    .io_connSS_35_data_qOutTask_bits(stealNet_io_connSS_35_data_qOutTask_bits),
    .io_connSS_36_ctrl_serveStealReq_ready(stealNet_io_connSS_36_ctrl_serveStealReq_ready),
    .io_connSS_36_ctrl_serveStealReq_valid(stealNet_io_connSS_36_ctrl_serveStealReq_valid),
    .io_connSS_36_ctrl_stealReq_ready(stealNet_io_connSS_36_ctrl_stealReq_ready),
    .io_connSS_36_ctrl_stealReq_valid(stealNet_io_connSS_36_ctrl_stealReq_valid),
    .io_connSS_36_data_availableTask_ready(stealNet_io_connSS_36_data_availableTask_ready),
    .io_connSS_36_data_availableTask_valid(stealNet_io_connSS_36_data_availableTask_valid),
    .io_connSS_36_data_availableTask_bits(stealNet_io_connSS_36_data_availableTask_bits),
    .io_connSS_36_data_qOutTask_ready(stealNet_io_connSS_36_data_qOutTask_ready),
    .io_connSS_36_data_qOutTask_valid(stealNet_io_connSS_36_data_qOutTask_valid),
    .io_connSS_36_data_qOutTask_bits(stealNet_io_connSS_36_data_qOutTask_bits),
    .io_connSS_37_ctrl_serveStealReq_ready(stealNet_io_connSS_37_ctrl_serveStealReq_ready),
    .io_connSS_37_ctrl_serveStealReq_valid(stealNet_io_connSS_37_ctrl_serveStealReq_valid),
    .io_connSS_37_ctrl_stealReq_ready(stealNet_io_connSS_37_ctrl_stealReq_ready),
    .io_connSS_37_ctrl_stealReq_valid(stealNet_io_connSS_37_ctrl_stealReq_valid),
    .io_connSS_37_data_availableTask_ready(stealNet_io_connSS_37_data_availableTask_ready),
    .io_connSS_37_data_availableTask_valid(stealNet_io_connSS_37_data_availableTask_valid),
    .io_connSS_37_data_availableTask_bits(stealNet_io_connSS_37_data_availableTask_bits),
    .io_connSS_37_data_qOutTask_ready(stealNet_io_connSS_37_data_qOutTask_ready),
    .io_connSS_37_data_qOutTask_valid(stealNet_io_connSS_37_data_qOutTask_valid),
    .io_connSS_37_data_qOutTask_bits(stealNet_io_connSS_37_data_qOutTask_bits),
    .io_connSS_38_ctrl_serveStealReq_ready(stealNet_io_connSS_38_ctrl_serveStealReq_ready),
    .io_connSS_38_ctrl_serveStealReq_valid(stealNet_io_connSS_38_ctrl_serveStealReq_valid),
    .io_connSS_38_ctrl_stealReq_ready(stealNet_io_connSS_38_ctrl_stealReq_ready),
    .io_connSS_38_ctrl_stealReq_valid(stealNet_io_connSS_38_ctrl_stealReq_valid),
    .io_connSS_38_data_availableTask_ready(stealNet_io_connSS_38_data_availableTask_ready),
    .io_connSS_38_data_availableTask_valid(stealNet_io_connSS_38_data_availableTask_valid),
    .io_connSS_38_data_availableTask_bits(stealNet_io_connSS_38_data_availableTask_bits),
    .io_connSS_38_data_qOutTask_ready(stealNet_io_connSS_38_data_qOutTask_ready),
    .io_connSS_38_data_qOutTask_valid(stealNet_io_connSS_38_data_qOutTask_valid),
    .io_connSS_38_data_qOutTask_bits(stealNet_io_connSS_38_data_qOutTask_bits),
    .io_connSS_39_ctrl_serveStealReq_ready(stealNet_io_connSS_39_ctrl_serveStealReq_ready),
    .io_connSS_39_ctrl_serveStealReq_valid(stealNet_io_connSS_39_ctrl_serveStealReq_valid),
    .io_connSS_39_ctrl_stealReq_ready(stealNet_io_connSS_39_ctrl_stealReq_ready),
    .io_connSS_39_ctrl_stealReq_valid(stealNet_io_connSS_39_ctrl_stealReq_valid),
    .io_connSS_39_data_availableTask_ready(stealNet_io_connSS_39_data_availableTask_ready),
    .io_connSS_39_data_availableTask_valid(stealNet_io_connSS_39_data_availableTask_valid),
    .io_connSS_39_data_availableTask_bits(stealNet_io_connSS_39_data_availableTask_bits),
    .io_connSS_39_data_qOutTask_ready(stealNet_io_connSS_39_data_qOutTask_ready),
    .io_connSS_39_data_qOutTask_valid(stealNet_io_connSS_39_data_qOutTask_valid),
    .io_connSS_39_data_qOutTask_bits(stealNet_io_connSS_39_data_qOutTask_bits),
    .io_connSS_40_ctrl_serveStealReq_ready(stealNet_io_connSS_40_ctrl_serveStealReq_ready),
    .io_connSS_40_ctrl_serveStealReq_valid(stealNet_io_connSS_40_ctrl_serveStealReq_valid),
    .io_connSS_40_ctrl_stealReq_ready(stealNet_io_connSS_40_ctrl_stealReq_ready),
    .io_connSS_40_ctrl_stealReq_valid(stealNet_io_connSS_40_ctrl_stealReq_valid),
    .io_connSS_40_data_availableTask_ready(stealNet_io_connSS_40_data_availableTask_ready),
    .io_connSS_40_data_availableTask_valid(stealNet_io_connSS_40_data_availableTask_valid),
    .io_connSS_40_data_availableTask_bits(stealNet_io_connSS_40_data_availableTask_bits),
    .io_connSS_40_data_qOutTask_ready(stealNet_io_connSS_40_data_qOutTask_ready),
    .io_connSS_40_data_qOutTask_valid(stealNet_io_connSS_40_data_qOutTask_valid),
    .io_connSS_40_data_qOutTask_bits(stealNet_io_connSS_40_data_qOutTask_bits),
    .io_connSS_41_ctrl_serveStealReq_ready(stealNet_io_connSS_41_ctrl_serveStealReq_ready),
    .io_connSS_41_ctrl_serveStealReq_valid(stealNet_io_connSS_41_ctrl_serveStealReq_valid),
    .io_connSS_41_ctrl_stealReq_ready(stealNet_io_connSS_41_ctrl_stealReq_ready),
    .io_connSS_41_ctrl_stealReq_valid(stealNet_io_connSS_41_ctrl_stealReq_valid),
    .io_connSS_41_data_availableTask_ready(stealNet_io_connSS_41_data_availableTask_ready),
    .io_connSS_41_data_availableTask_valid(stealNet_io_connSS_41_data_availableTask_valid),
    .io_connSS_41_data_availableTask_bits(stealNet_io_connSS_41_data_availableTask_bits),
    .io_connSS_41_data_qOutTask_ready(stealNet_io_connSS_41_data_qOutTask_ready),
    .io_connSS_41_data_qOutTask_valid(stealNet_io_connSS_41_data_qOutTask_valid),
    .io_connSS_41_data_qOutTask_bits(stealNet_io_connSS_41_data_qOutTask_bits),
    .io_connSS_42_ctrl_serveStealReq_ready(stealNet_io_connSS_42_ctrl_serveStealReq_ready),
    .io_connSS_42_ctrl_serveStealReq_valid(stealNet_io_connSS_42_ctrl_serveStealReq_valid),
    .io_connSS_42_ctrl_stealReq_ready(stealNet_io_connSS_42_ctrl_stealReq_ready),
    .io_connSS_42_ctrl_stealReq_valid(stealNet_io_connSS_42_ctrl_stealReq_valid),
    .io_connSS_42_data_availableTask_ready(stealNet_io_connSS_42_data_availableTask_ready),
    .io_connSS_42_data_availableTask_valid(stealNet_io_connSS_42_data_availableTask_valid),
    .io_connSS_42_data_availableTask_bits(stealNet_io_connSS_42_data_availableTask_bits),
    .io_connSS_42_data_qOutTask_ready(stealNet_io_connSS_42_data_qOutTask_ready),
    .io_connSS_42_data_qOutTask_valid(stealNet_io_connSS_42_data_qOutTask_valid),
    .io_connSS_42_data_qOutTask_bits(stealNet_io_connSS_42_data_qOutTask_bits),
    .io_connSS_43_ctrl_serveStealReq_ready(stealNet_io_connSS_43_ctrl_serveStealReq_ready),
    .io_connSS_43_ctrl_serveStealReq_valid(stealNet_io_connSS_43_ctrl_serveStealReq_valid),
    .io_connSS_43_ctrl_stealReq_ready(stealNet_io_connSS_43_ctrl_stealReq_ready),
    .io_connSS_43_ctrl_stealReq_valid(stealNet_io_connSS_43_ctrl_stealReq_valid),
    .io_connSS_43_data_availableTask_ready(stealNet_io_connSS_43_data_availableTask_ready),
    .io_connSS_43_data_availableTask_valid(stealNet_io_connSS_43_data_availableTask_valid),
    .io_connSS_43_data_availableTask_bits(stealNet_io_connSS_43_data_availableTask_bits),
    .io_connSS_43_data_qOutTask_ready(stealNet_io_connSS_43_data_qOutTask_ready),
    .io_connSS_43_data_qOutTask_valid(stealNet_io_connSS_43_data_qOutTask_valid),
    .io_connSS_43_data_qOutTask_bits(stealNet_io_connSS_43_data_qOutTask_bits),
    .io_connSS_44_ctrl_serveStealReq_ready(stealNet_io_connSS_44_ctrl_serveStealReq_ready),
    .io_connSS_44_ctrl_serveStealReq_valid(stealNet_io_connSS_44_ctrl_serveStealReq_valid),
    .io_connSS_44_ctrl_stealReq_ready(stealNet_io_connSS_44_ctrl_stealReq_ready),
    .io_connSS_44_ctrl_stealReq_valid(stealNet_io_connSS_44_ctrl_stealReq_valid),
    .io_connSS_44_data_availableTask_ready(stealNet_io_connSS_44_data_availableTask_ready),
    .io_connSS_44_data_availableTask_valid(stealNet_io_connSS_44_data_availableTask_valid),
    .io_connSS_44_data_availableTask_bits(stealNet_io_connSS_44_data_availableTask_bits),
    .io_connSS_44_data_qOutTask_ready(stealNet_io_connSS_44_data_qOutTask_ready),
    .io_connSS_44_data_qOutTask_valid(stealNet_io_connSS_44_data_qOutTask_valid),
    .io_connSS_44_data_qOutTask_bits(stealNet_io_connSS_44_data_qOutTask_bits),
    .io_connSS_45_ctrl_serveStealReq_ready(stealNet_io_connSS_45_ctrl_serveStealReq_ready),
    .io_connSS_45_ctrl_serveStealReq_valid(stealNet_io_connSS_45_ctrl_serveStealReq_valid),
    .io_connSS_45_ctrl_stealReq_ready(stealNet_io_connSS_45_ctrl_stealReq_ready),
    .io_connSS_45_ctrl_stealReq_valid(stealNet_io_connSS_45_ctrl_stealReq_valid),
    .io_connSS_45_data_availableTask_ready(stealNet_io_connSS_45_data_availableTask_ready),
    .io_connSS_45_data_availableTask_valid(stealNet_io_connSS_45_data_availableTask_valid),
    .io_connSS_45_data_availableTask_bits(stealNet_io_connSS_45_data_availableTask_bits),
    .io_connSS_45_data_qOutTask_ready(stealNet_io_connSS_45_data_qOutTask_ready),
    .io_connSS_45_data_qOutTask_valid(stealNet_io_connSS_45_data_qOutTask_valid),
    .io_connSS_45_data_qOutTask_bits(stealNet_io_connSS_45_data_qOutTask_bits),
    .io_connSS_46_ctrl_serveStealReq_ready(stealNet_io_connSS_46_ctrl_serveStealReq_ready),
    .io_connSS_46_ctrl_serveStealReq_valid(stealNet_io_connSS_46_ctrl_serveStealReq_valid),
    .io_connSS_46_ctrl_stealReq_ready(stealNet_io_connSS_46_ctrl_stealReq_ready),
    .io_connSS_46_ctrl_stealReq_valid(stealNet_io_connSS_46_ctrl_stealReq_valid),
    .io_connSS_46_data_availableTask_ready(stealNet_io_connSS_46_data_availableTask_ready),
    .io_connSS_46_data_availableTask_valid(stealNet_io_connSS_46_data_availableTask_valid),
    .io_connSS_46_data_availableTask_bits(stealNet_io_connSS_46_data_availableTask_bits),
    .io_connSS_46_data_qOutTask_ready(stealNet_io_connSS_46_data_qOutTask_ready),
    .io_connSS_46_data_qOutTask_valid(stealNet_io_connSS_46_data_qOutTask_valid),
    .io_connSS_46_data_qOutTask_bits(stealNet_io_connSS_46_data_qOutTask_bits),
    .io_connSS_47_ctrl_serveStealReq_ready(stealNet_io_connSS_47_ctrl_serveStealReq_ready),
    .io_connSS_47_ctrl_serveStealReq_valid(stealNet_io_connSS_47_ctrl_serveStealReq_valid),
    .io_connSS_47_ctrl_stealReq_ready(stealNet_io_connSS_47_ctrl_stealReq_ready),
    .io_connSS_47_ctrl_stealReq_valid(stealNet_io_connSS_47_ctrl_stealReq_valid),
    .io_connSS_47_data_availableTask_ready(stealNet_io_connSS_47_data_availableTask_ready),
    .io_connSS_47_data_availableTask_valid(stealNet_io_connSS_47_data_availableTask_valid),
    .io_connSS_47_data_availableTask_bits(stealNet_io_connSS_47_data_availableTask_bits),
    .io_connSS_47_data_qOutTask_ready(stealNet_io_connSS_47_data_qOutTask_ready),
    .io_connSS_47_data_qOutTask_valid(stealNet_io_connSS_47_data_qOutTask_valid),
    .io_connSS_47_data_qOutTask_bits(stealNet_io_connSS_47_data_qOutTask_bits),
    .io_connSS_48_ctrl_serveStealReq_ready(stealNet_io_connSS_48_ctrl_serveStealReq_ready),
    .io_connSS_48_ctrl_serveStealReq_valid(stealNet_io_connSS_48_ctrl_serveStealReq_valid),
    .io_connSS_48_ctrl_stealReq_ready(stealNet_io_connSS_48_ctrl_stealReq_ready),
    .io_connSS_48_ctrl_stealReq_valid(stealNet_io_connSS_48_ctrl_stealReq_valid),
    .io_connSS_48_data_availableTask_ready(stealNet_io_connSS_48_data_availableTask_ready),
    .io_connSS_48_data_availableTask_valid(stealNet_io_connSS_48_data_availableTask_valid),
    .io_connSS_48_data_availableTask_bits(stealNet_io_connSS_48_data_availableTask_bits),
    .io_connSS_48_data_qOutTask_ready(stealNet_io_connSS_48_data_qOutTask_ready),
    .io_connSS_48_data_qOutTask_valid(stealNet_io_connSS_48_data_qOutTask_valid),
    .io_connSS_48_data_qOutTask_bits(stealNet_io_connSS_48_data_qOutTask_bits),
    .io_connSS_49_ctrl_serveStealReq_ready(stealNet_io_connSS_49_ctrl_serveStealReq_ready),
    .io_connSS_49_ctrl_serveStealReq_valid(stealNet_io_connSS_49_ctrl_serveStealReq_valid),
    .io_connSS_49_ctrl_stealReq_ready(stealNet_io_connSS_49_ctrl_stealReq_ready),
    .io_connSS_49_ctrl_stealReq_valid(stealNet_io_connSS_49_ctrl_stealReq_valid),
    .io_connSS_49_data_availableTask_ready(stealNet_io_connSS_49_data_availableTask_ready),
    .io_connSS_49_data_availableTask_valid(stealNet_io_connSS_49_data_availableTask_valid),
    .io_connSS_49_data_availableTask_bits(stealNet_io_connSS_49_data_availableTask_bits),
    .io_connSS_49_data_qOutTask_ready(stealNet_io_connSS_49_data_qOutTask_ready),
    .io_connSS_49_data_qOutTask_valid(stealNet_io_connSS_49_data_qOutTask_valid),
    .io_connSS_49_data_qOutTask_bits(stealNet_io_connSS_49_data_qOutTask_bits),
    .io_connSS_50_ctrl_serveStealReq_ready(stealNet_io_connSS_50_ctrl_serveStealReq_ready),
    .io_connSS_50_ctrl_serveStealReq_valid(stealNet_io_connSS_50_ctrl_serveStealReq_valid),
    .io_connSS_50_ctrl_stealReq_ready(stealNet_io_connSS_50_ctrl_stealReq_ready),
    .io_connSS_50_ctrl_stealReq_valid(stealNet_io_connSS_50_ctrl_stealReq_valid),
    .io_connSS_50_data_availableTask_ready(stealNet_io_connSS_50_data_availableTask_ready),
    .io_connSS_50_data_availableTask_valid(stealNet_io_connSS_50_data_availableTask_valid),
    .io_connSS_50_data_availableTask_bits(stealNet_io_connSS_50_data_availableTask_bits),
    .io_connSS_50_data_qOutTask_ready(stealNet_io_connSS_50_data_qOutTask_ready),
    .io_connSS_50_data_qOutTask_valid(stealNet_io_connSS_50_data_qOutTask_valid),
    .io_connSS_50_data_qOutTask_bits(stealNet_io_connSS_50_data_qOutTask_bits),
    .io_connSS_51_ctrl_serveStealReq_ready(stealNet_io_connSS_51_ctrl_serveStealReq_ready),
    .io_connSS_51_ctrl_serveStealReq_valid(stealNet_io_connSS_51_ctrl_serveStealReq_valid),
    .io_connSS_51_ctrl_stealReq_ready(stealNet_io_connSS_51_ctrl_stealReq_ready),
    .io_connSS_51_ctrl_stealReq_valid(stealNet_io_connSS_51_ctrl_stealReq_valid),
    .io_connSS_51_data_availableTask_ready(stealNet_io_connSS_51_data_availableTask_ready),
    .io_connSS_51_data_availableTask_valid(stealNet_io_connSS_51_data_availableTask_valid),
    .io_connSS_51_data_availableTask_bits(stealNet_io_connSS_51_data_availableTask_bits),
    .io_connSS_51_data_qOutTask_ready(stealNet_io_connSS_51_data_qOutTask_ready),
    .io_connSS_51_data_qOutTask_valid(stealNet_io_connSS_51_data_qOutTask_valid),
    .io_connSS_51_data_qOutTask_bits(stealNet_io_connSS_51_data_qOutTask_bits),
    .io_connSS_52_ctrl_serveStealReq_ready(stealNet_io_connSS_52_ctrl_serveStealReq_ready),
    .io_connSS_52_ctrl_serveStealReq_valid(stealNet_io_connSS_52_ctrl_serveStealReq_valid),
    .io_connSS_52_ctrl_stealReq_ready(stealNet_io_connSS_52_ctrl_stealReq_ready),
    .io_connSS_52_ctrl_stealReq_valid(stealNet_io_connSS_52_ctrl_stealReq_valid),
    .io_connSS_52_data_availableTask_ready(stealNet_io_connSS_52_data_availableTask_ready),
    .io_connSS_52_data_availableTask_valid(stealNet_io_connSS_52_data_availableTask_valid),
    .io_connSS_52_data_availableTask_bits(stealNet_io_connSS_52_data_availableTask_bits),
    .io_connSS_52_data_qOutTask_ready(stealNet_io_connSS_52_data_qOutTask_ready),
    .io_connSS_52_data_qOutTask_valid(stealNet_io_connSS_52_data_qOutTask_valid),
    .io_connSS_52_data_qOutTask_bits(stealNet_io_connSS_52_data_qOutTask_bits),
    .io_connSS_53_ctrl_serveStealReq_ready(stealNet_io_connSS_53_ctrl_serveStealReq_ready),
    .io_connSS_53_ctrl_serveStealReq_valid(stealNet_io_connSS_53_ctrl_serveStealReq_valid),
    .io_connSS_53_ctrl_stealReq_ready(stealNet_io_connSS_53_ctrl_stealReq_ready),
    .io_connSS_53_ctrl_stealReq_valid(stealNet_io_connSS_53_ctrl_stealReq_valid),
    .io_connSS_53_data_availableTask_ready(stealNet_io_connSS_53_data_availableTask_ready),
    .io_connSS_53_data_availableTask_valid(stealNet_io_connSS_53_data_availableTask_valid),
    .io_connSS_53_data_availableTask_bits(stealNet_io_connSS_53_data_availableTask_bits),
    .io_connSS_53_data_qOutTask_ready(stealNet_io_connSS_53_data_qOutTask_ready),
    .io_connSS_53_data_qOutTask_valid(stealNet_io_connSS_53_data_qOutTask_valid),
    .io_connSS_53_data_qOutTask_bits(stealNet_io_connSS_53_data_qOutTask_bits),
    .io_connSS_54_ctrl_serveStealReq_ready(stealNet_io_connSS_54_ctrl_serveStealReq_ready),
    .io_connSS_54_ctrl_serveStealReq_valid(stealNet_io_connSS_54_ctrl_serveStealReq_valid),
    .io_connSS_54_ctrl_stealReq_ready(stealNet_io_connSS_54_ctrl_stealReq_ready),
    .io_connSS_54_ctrl_stealReq_valid(stealNet_io_connSS_54_ctrl_stealReq_valid),
    .io_connSS_54_data_availableTask_ready(stealNet_io_connSS_54_data_availableTask_ready),
    .io_connSS_54_data_availableTask_valid(stealNet_io_connSS_54_data_availableTask_valid),
    .io_connSS_54_data_availableTask_bits(stealNet_io_connSS_54_data_availableTask_bits),
    .io_connSS_54_data_qOutTask_ready(stealNet_io_connSS_54_data_qOutTask_ready),
    .io_connSS_54_data_qOutTask_valid(stealNet_io_connSS_54_data_qOutTask_valid),
    .io_connSS_54_data_qOutTask_bits(stealNet_io_connSS_54_data_qOutTask_bits),
    .io_connSS_55_ctrl_serveStealReq_ready(stealNet_io_connSS_55_ctrl_serveStealReq_ready),
    .io_connSS_55_ctrl_serveStealReq_valid(stealNet_io_connSS_55_ctrl_serveStealReq_valid),
    .io_connSS_55_ctrl_stealReq_ready(stealNet_io_connSS_55_ctrl_stealReq_ready),
    .io_connSS_55_ctrl_stealReq_valid(stealNet_io_connSS_55_ctrl_stealReq_valid),
    .io_connSS_55_data_availableTask_ready(stealNet_io_connSS_55_data_availableTask_ready),
    .io_connSS_55_data_availableTask_valid(stealNet_io_connSS_55_data_availableTask_valid),
    .io_connSS_55_data_availableTask_bits(stealNet_io_connSS_55_data_availableTask_bits),
    .io_connSS_55_data_qOutTask_ready(stealNet_io_connSS_55_data_qOutTask_ready),
    .io_connSS_55_data_qOutTask_valid(stealNet_io_connSS_55_data_qOutTask_valid),
    .io_connSS_55_data_qOutTask_bits(stealNet_io_connSS_55_data_qOutTask_bits),
    .io_connSS_56_ctrl_serveStealReq_ready(stealNet_io_connSS_56_ctrl_serveStealReq_ready),
    .io_connSS_56_ctrl_serveStealReq_valid(stealNet_io_connSS_56_ctrl_serveStealReq_valid),
    .io_connSS_56_ctrl_stealReq_ready(stealNet_io_connSS_56_ctrl_stealReq_ready),
    .io_connSS_56_ctrl_stealReq_valid(stealNet_io_connSS_56_ctrl_stealReq_valid),
    .io_connSS_56_data_availableTask_ready(stealNet_io_connSS_56_data_availableTask_ready),
    .io_connSS_56_data_availableTask_valid(stealNet_io_connSS_56_data_availableTask_valid),
    .io_connSS_56_data_availableTask_bits(stealNet_io_connSS_56_data_availableTask_bits),
    .io_connSS_56_data_qOutTask_ready(stealNet_io_connSS_56_data_qOutTask_ready),
    .io_connSS_56_data_qOutTask_valid(stealNet_io_connSS_56_data_qOutTask_valid),
    .io_connSS_56_data_qOutTask_bits(stealNet_io_connSS_56_data_qOutTask_bits),
    .io_connSS_57_ctrl_serveStealReq_ready(stealNet_io_connSS_57_ctrl_serveStealReq_ready),
    .io_connSS_57_ctrl_serveStealReq_valid(stealNet_io_connSS_57_ctrl_serveStealReq_valid),
    .io_connSS_57_ctrl_stealReq_ready(stealNet_io_connSS_57_ctrl_stealReq_ready),
    .io_connSS_57_ctrl_stealReq_valid(stealNet_io_connSS_57_ctrl_stealReq_valid),
    .io_connSS_57_data_availableTask_ready(stealNet_io_connSS_57_data_availableTask_ready),
    .io_connSS_57_data_availableTask_valid(stealNet_io_connSS_57_data_availableTask_valid),
    .io_connSS_57_data_availableTask_bits(stealNet_io_connSS_57_data_availableTask_bits),
    .io_connSS_57_data_qOutTask_ready(stealNet_io_connSS_57_data_qOutTask_ready),
    .io_connSS_57_data_qOutTask_valid(stealNet_io_connSS_57_data_qOutTask_valid),
    .io_connSS_57_data_qOutTask_bits(stealNet_io_connSS_57_data_qOutTask_bits),
    .io_connSS_58_ctrl_serveStealReq_ready(stealNet_io_connSS_58_ctrl_serveStealReq_ready),
    .io_connSS_58_ctrl_serveStealReq_valid(stealNet_io_connSS_58_ctrl_serveStealReq_valid),
    .io_connSS_58_ctrl_stealReq_ready(stealNet_io_connSS_58_ctrl_stealReq_ready),
    .io_connSS_58_ctrl_stealReq_valid(stealNet_io_connSS_58_ctrl_stealReq_valid),
    .io_connSS_58_data_availableTask_ready(stealNet_io_connSS_58_data_availableTask_ready),
    .io_connSS_58_data_availableTask_valid(stealNet_io_connSS_58_data_availableTask_valid),
    .io_connSS_58_data_availableTask_bits(stealNet_io_connSS_58_data_availableTask_bits),
    .io_connSS_58_data_qOutTask_ready(stealNet_io_connSS_58_data_qOutTask_ready),
    .io_connSS_58_data_qOutTask_valid(stealNet_io_connSS_58_data_qOutTask_valid),
    .io_connSS_58_data_qOutTask_bits(stealNet_io_connSS_58_data_qOutTask_bits),
    .io_connSS_59_ctrl_serveStealReq_ready(stealNet_io_connSS_59_ctrl_serveStealReq_ready),
    .io_connSS_59_ctrl_serveStealReq_valid(stealNet_io_connSS_59_ctrl_serveStealReq_valid),
    .io_connSS_59_ctrl_stealReq_ready(stealNet_io_connSS_59_ctrl_stealReq_ready),
    .io_connSS_59_ctrl_stealReq_valid(stealNet_io_connSS_59_ctrl_stealReq_valid),
    .io_connSS_59_data_availableTask_ready(stealNet_io_connSS_59_data_availableTask_ready),
    .io_connSS_59_data_availableTask_valid(stealNet_io_connSS_59_data_availableTask_valid),
    .io_connSS_59_data_availableTask_bits(stealNet_io_connSS_59_data_availableTask_bits),
    .io_connSS_59_data_qOutTask_ready(stealNet_io_connSS_59_data_qOutTask_ready),
    .io_connSS_59_data_qOutTask_valid(stealNet_io_connSS_59_data_qOutTask_valid),
    .io_connSS_59_data_qOutTask_bits(stealNet_io_connSS_59_data_qOutTask_bits),
    .io_connSS_60_ctrl_serveStealReq_ready(stealNet_io_connSS_60_ctrl_serveStealReq_ready),
    .io_connSS_60_ctrl_serveStealReq_valid(stealNet_io_connSS_60_ctrl_serveStealReq_valid),
    .io_connSS_60_ctrl_stealReq_ready(stealNet_io_connSS_60_ctrl_stealReq_ready),
    .io_connSS_60_ctrl_stealReq_valid(stealNet_io_connSS_60_ctrl_stealReq_valid),
    .io_connSS_60_data_availableTask_ready(stealNet_io_connSS_60_data_availableTask_ready),
    .io_connSS_60_data_availableTask_valid(stealNet_io_connSS_60_data_availableTask_valid),
    .io_connSS_60_data_availableTask_bits(stealNet_io_connSS_60_data_availableTask_bits),
    .io_connSS_60_data_qOutTask_ready(stealNet_io_connSS_60_data_qOutTask_ready),
    .io_connSS_60_data_qOutTask_valid(stealNet_io_connSS_60_data_qOutTask_valid),
    .io_connSS_60_data_qOutTask_bits(stealNet_io_connSS_60_data_qOutTask_bits),
    .io_connSS_61_ctrl_serveStealReq_ready(stealNet_io_connSS_61_ctrl_serveStealReq_ready),
    .io_connSS_61_ctrl_serveStealReq_valid(stealNet_io_connSS_61_ctrl_serveStealReq_valid),
    .io_connSS_61_ctrl_stealReq_ready(stealNet_io_connSS_61_ctrl_stealReq_ready),
    .io_connSS_61_ctrl_stealReq_valid(stealNet_io_connSS_61_ctrl_stealReq_valid),
    .io_connSS_61_data_availableTask_ready(stealNet_io_connSS_61_data_availableTask_ready),
    .io_connSS_61_data_availableTask_valid(stealNet_io_connSS_61_data_availableTask_valid),
    .io_connSS_61_data_availableTask_bits(stealNet_io_connSS_61_data_availableTask_bits),
    .io_connSS_61_data_qOutTask_ready(stealNet_io_connSS_61_data_qOutTask_ready),
    .io_connSS_61_data_qOutTask_valid(stealNet_io_connSS_61_data_qOutTask_valid),
    .io_connSS_61_data_qOutTask_bits(stealNet_io_connSS_61_data_qOutTask_bits),
    .io_connSS_62_ctrl_serveStealReq_ready(stealNet_io_connSS_62_ctrl_serveStealReq_ready),
    .io_connSS_62_ctrl_serveStealReq_valid(stealNet_io_connSS_62_ctrl_serveStealReq_valid),
    .io_connSS_62_ctrl_stealReq_ready(stealNet_io_connSS_62_ctrl_stealReq_ready),
    .io_connSS_62_ctrl_stealReq_valid(stealNet_io_connSS_62_ctrl_stealReq_valid),
    .io_connSS_62_data_availableTask_ready(stealNet_io_connSS_62_data_availableTask_ready),
    .io_connSS_62_data_availableTask_valid(stealNet_io_connSS_62_data_availableTask_valid),
    .io_connSS_62_data_availableTask_bits(stealNet_io_connSS_62_data_availableTask_bits),
    .io_connSS_62_data_qOutTask_ready(stealNet_io_connSS_62_data_qOutTask_ready),
    .io_connSS_62_data_qOutTask_valid(stealNet_io_connSS_62_data_qOutTask_valid),
    .io_connSS_62_data_qOutTask_bits(stealNet_io_connSS_62_data_qOutTask_bits),
    .io_connSS_63_ctrl_serveStealReq_ready(stealNet_io_connSS_63_ctrl_serveStealReq_ready),
    .io_connSS_63_ctrl_serveStealReq_valid(stealNet_io_connSS_63_ctrl_serveStealReq_valid),
    .io_connSS_63_ctrl_stealReq_ready(stealNet_io_connSS_63_ctrl_stealReq_ready),
    .io_connSS_63_ctrl_stealReq_valid(stealNet_io_connSS_63_ctrl_stealReq_valid),
    .io_connSS_63_data_availableTask_ready(stealNet_io_connSS_63_data_availableTask_ready),
    .io_connSS_63_data_availableTask_valid(stealNet_io_connSS_63_data_availableTask_valid),
    .io_connSS_63_data_availableTask_bits(stealNet_io_connSS_63_data_availableTask_bits),
    .io_connSS_63_data_qOutTask_ready(stealNet_io_connSS_63_data_qOutTask_ready),
    .io_connSS_63_data_qOutTask_valid(stealNet_io_connSS_63_data_qOutTask_valid),
    .io_connSS_63_data_qOutTask_bits(stealNet_io_connSS_63_data_qOutTask_bits),
    .io_connSS_64_ctrl_serveStealReq_ready(stealNet_io_connSS_64_ctrl_serveStealReq_ready),
    .io_connSS_64_ctrl_serveStealReq_valid(stealNet_io_connSS_64_ctrl_serveStealReq_valid),
    .io_connSS_64_ctrl_stealReq_ready(stealNet_io_connSS_64_ctrl_stealReq_ready),
    .io_connSS_64_ctrl_stealReq_valid(stealNet_io_connSS_64_ctrl_stealReq_valid),
    .io_connSS_64_data_availableTask_ready(stealNet_io_connSS_64_data_availableTask_ready),
    .io_connSS_64_data_availableTask_valid(stealNet_io_connSS_64_data_availableTask_valid),
    .io_connSS_64_data_availableTask_bits(stealNet_io_connSS_64_data_availableTask_bits),
    .io_connSS_64_data_qOutTask_ready(stealNet_io_connSS_64_data_qOutTask_ready),
    .io_connSS_64_data_qOutTask_valid(stealNet_io_connSS_64_data_qOutTask_valid),
    .io_connSS_64_data_qOutTask_bits(stealNet_io_connSS_64_data_qOutTask_bits),
    .io_connSS_65_ctrl_serveStealReq_ready(stealNet_io_connSS_65_ctrl_serveStealReq_ready),
    .io_connSS_65_ctrl_serveStealReq_valid(stealNet_io_connSS_65_ctrl_serveStealReq_valid),
    .io_connSS_65_ctrl_stealReq_ready(stealNet_io_connSS_65_ctrl_stealReq_ready),
    .io_connSS_65_ctrl_stealReq_valid(stealNet_io_connSS_65_ctrl_stealReq_valid),
    .io_connSS_65_data_availableTask_ready(stealNet_io_connSS_65_data_availableTask_ready),
    .io_connSS_65_data_availableTask_valid(stealNet_io_connSS_65_data_availableTask_valid),
    .io_connSS_65_data_availableTask_bits(stealNet_io_connSS_65_data_availableTask_bits),
    .io_connSS_65_data_qOutTask_ready(stealNet_io_connSS_65_data_qOutTask_ready),
    .io_connSS_65_data_qOutTask_valid(stealNet_io_connSS_65_data_qOutTask_valid),
    .io_connSS_65_data_qOutTask_bits(stealNet_io_connSS_65_data_qOutTask_bits),
    .io_connSS_66_ctrl_serveStealReq_ready(stealNet_io_connSS_66_ctrl_serveStealReq_ready),
    .io_connSS_66_ctrl_serveStealReq_valid(stealNet_io_connSS_66_ctrl_serveStealReq_valid),
    .io_connSS_66_ctrl_stealReq_ready(stealNet_io_connSS_66_ctrl_stealReq_ready),
    .io_connSS_66_ctrl_stealReq_valid(stealNet_io_connSS_66_ctrl_stealReq_valid),
    .io_connSS_66_data_availableTask_ready(stealNet_io_connSS_66_data_availableTask_ready),
    .io_connSS_66_data_availableTask_valid(stealNet_io_connSS_66_data_availableTask_valid),
    .io_connSS_66_data_availableTask_bits(stealNet_io_connSS_66_data_availableTask_bits),
    .io_connSS_66_data_qOutTask_ready(stealNet_io_connSS_66_data_qOutTask_ready),
    .io_connSS_66_data_qOutTask_valid(stealNet_io_connSS_66_data_qOutTask_valid),
    .io_connSS_66_data_qOutTask_bits(stealNet_io_connSS_66_data_qOutTask_bits),
    .io_ntwDataUnitOccupancyVSS_0(stealNet_io_ntwDataUnitOccupancyVSS_0)
  );
  stealServer stealServers_0 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_0_clock),
    .reset(stealServers_0_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_0_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_0_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_0_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_0_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_0_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_0_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_0_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_0_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_0_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_0_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_0_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_0_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_0_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_0_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_0_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_0_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_0_io_connQ_pop_bits)
  );
  stealServer stealServers_1 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_1_clock),
    .reset(stealServers_1_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_1_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_1_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_1_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_1_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_1_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_1_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_1_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_1_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_1_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_1_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_1_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_1_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_1_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_1_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_1_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_1_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_1_io_connQ_pop_bits)
  );
  stealServer stealServers_2 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_2_clock),
    .reset(stealServers_2_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_2_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_2_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_2_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_2_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_2_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_2_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_2_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_2_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_2_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_2_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_2_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_2_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_2_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_2_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_2_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_2_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_2_io_connQ_pop_bits)
  );
  stealServer stealServers_3 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_3_clock),
    .reset(stealServers_3_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_3_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_3_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_3_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_3_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_3_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_3_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_3_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_3_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_3_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_3_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_3_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_3_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_3_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_3_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_3_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_3_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_3_io_connQ_pop_bits)
  );
  stealServer stealServers_4 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_4_clock),
    .reset(stealServers_4_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_4_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_4_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_4_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_4_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_4_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_4_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_4_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_4_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_4_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_4_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_4_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_4_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_4_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_4_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_4_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_4_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_4_io_connQ_pop_bits)
  );
  stealServer stealServers_5 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_5_clock),
    .reset(stealServers_5_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_5_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_5_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_5_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_5_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_5_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_5_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_5_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_5_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_5_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_5_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_5_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_5_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_5_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_5_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_5_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_5_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_5_io_connQ_pop_bits)
  );
  stealServer stealServers_6 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_6_clock),
    .reset(stealServers_6_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_6_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_6_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_6_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_6_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_6_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_6_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_6_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_6_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_6_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_6_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_6_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_6_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_6_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_6_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_6_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_6_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_6_io_connQ_pop_bits)
  );
  stealServer stealServers_7 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_7_clock),
    .reset(stealServers_7_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_7_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_7_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_7_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_7_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_7_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_7_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_7_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_7_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_7_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_7_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_7_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_7_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_7_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_7_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_7_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_7_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_7_io_connQ_pop_bits)
  );
  stealServer stealServers_8 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_8_clock),
    .reset(stealServers_8_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_8_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_8_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_8_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_8_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_8_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_8_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_8_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_8_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_8_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_8_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_8_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_8_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_8_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_8_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_8_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_8_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_8_io_connQ_pop_bits)
  );
  stealServer stealServers_9 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_9_clock),
    .reset(stealServers_9_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_9_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_9_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_9_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_9_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_9_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_9_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_9_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_9_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_9_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_9_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_9_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_9_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_9_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_9_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_9_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_9_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_9_io_connQ_pop_bits)
  );
  stealServer stealServers_10 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_10_clock),
    .reset(stealServers_10_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_10_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_10_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_10_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_10_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_10_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_10_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_10_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_10_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_10_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_10_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_10_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_10_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_10_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_10_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_10_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_10_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_10_io_connQ_pop_bits)
  );
  stealServer stealServers_11 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_11_clock),
    .reset(stealServers_11_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_11_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_11_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_11_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_11_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_11_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_11_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_11_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_11_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_11_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_11_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_11_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_11_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_11_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_11_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_11_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_11_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_11_io_connQ_pop_bits)
  );
  stealServer stealServers_12 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_12_clock),
    .reset(stealServers_12_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_12_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_12_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_12_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_12_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_12_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_12_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_12_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_12_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_12_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_12_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_12_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_12_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_12_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_12_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_12_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_12_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_12_io_connQ_pop_bits)
  );
  stealServer stealServers_13 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_13_clock),
    .reset(stealServers_13_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_13_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_13_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_13_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_13_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_13_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_13_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_13_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_13_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_13_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_13_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_13_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_13_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_13_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_13_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_13_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_13_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_13_io_connQ_pop_bits)
  );
  stealServer stealServers_14 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_14_clock),
    .reset(stealServers_14_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_14_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_14_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_14_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_14_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_14_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_14_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_14_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_14_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_14_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_14_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_14_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_14_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_14_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_14_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_14_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_14_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_14_io_connQ_pop_bits)
  );
  stealServer stealServers_15 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_15_clock),
    .reset(stealServers_15_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_15_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_15_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_15_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_15_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_15_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_15_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_15_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_15_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_15_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_15_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_15_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_15_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_15_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_15_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_15_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_15_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_15_io_connQ_pop_bits)
  );
  stealServer stealServers_16 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_16_clock),
    .reset(stealServers_16_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_16_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_16_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_16_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_16_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_16_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_16_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_16_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_16_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_16_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_16_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_16_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_16_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_16_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_16_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_16_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_16_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_16_io_connQ_pop_bits)
  );
  stealServer stealServers_17 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_17_clock),
    .reset(stealServers_17_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_17_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_17_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_17_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_17_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_17_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_17_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_17_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_17_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_17_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_17_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_17_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_17_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_17_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_17_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_17_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_17_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_17_io_connQ_pop_bits)
  );
  stealServer stealServers_18 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_18_clock),
    .reset(stealServers_18_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_18_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_18_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_18_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_18_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_18_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_18_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_18_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_18_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_18_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_18_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_18_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_18_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_18_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_18_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_18_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_18_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_18_io_connQ_pop_bits)
  );
  stealServer stealServers_19 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_19_clock),
    .reset(stealServers_19_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_19_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_19_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_19_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_19_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_19_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_19_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_19_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_19_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_19_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_19_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_19_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_19_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_19_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_19_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_19_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_19_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_19_io_connQ_pop_bits)
  );
  stealServer stealServers_20 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_20_clock),
    .reset(stealServers_20_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_20_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_20_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_20_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_20_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_20_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_20_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_20_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_20_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_20_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_20_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_20_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_20_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_20_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_20_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_20_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_20_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_20_io_connQ_pop_bits)
  );
  stealServer stealServers_21 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_21_clock),
    .reset(stealServers_21_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_21_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_21_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_21_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_21_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_21_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_21_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_21_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_21_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_21_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_21_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_21_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_21_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_21_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_21_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_21_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_21_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_21_io_connQ_pop_bits)
  );
  stealServer stealServers_22 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_22_clock),
    .reset(stealServers_22_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_22_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_22_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_22_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_22_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_22_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_22_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_22_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_22_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_22_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_22_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_22_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_22_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_22_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_22_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_22_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_22_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_22_io_connQ_pop_bits)
  );
  stealServer stealServers_23 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_23_clock),
    .reset(stealServers_23_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_23_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_23_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_23_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_23_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_23_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_23_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_23_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_23_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_23_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_23_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_23_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_23_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_23_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_23_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_23_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_23_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_23_io_connQ_pop_bits)
  );
  stealServer stealServers_24 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_24_clock),
    .reset(stealServers_24_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_24_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_24_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_24_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_24_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_24_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_24_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_24_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_24_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_24_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_24_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_24_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_24_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_24_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_24_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_24_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_24_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_24_io_connQ_pop_bits)
  );
  stealServer stealServers_25 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_25_clock),
    .reset(stealServers_25_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_25_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_25_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_25_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_25_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_25_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_25_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_25_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_25_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_25_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_25_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_25_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_25_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_25_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_25_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_25_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_25_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_25_io_connQ_pop_bits)
  );
  stealServer stealServers_26 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_26_clock),
    .reset(stealServers_26_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_26_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_26_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_26_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_26_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_26_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_26_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_26_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_26_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_26_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_26_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_26_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_26_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_26_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_26_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_26_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_26_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_26_io_connQ_pop_bits)
  );
  stealServer stealServers_27 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_27_clock),
    .reset(stealServers_27_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_27_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_27_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_27_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_27_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_27_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_27_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_27_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_27_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_27_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_27_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_27_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_27_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_27_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_27_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_27_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_27_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_27_io_connQ_pop_bits)
  );
  stealServer stealServers_28 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_28_clock),
    .reset(stealServers_28_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_28_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_28_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_28_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_28_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_28_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_28_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_28_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_28_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_28_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_28_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_28_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_28_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_28_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_28_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_28_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_28_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_28_io_connQ_pop_bits)
  );
  stealServer stealServers_29 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_29_clock),
    .reset(stealServers_29_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_29_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_29_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_29_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_29_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_29_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_29_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_29_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_29_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_29_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_29_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_29_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_29_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_29_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_29_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_29_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_29_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_29_io_connQ_pop_bits)
  );
  stealServer stealServers_30 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_30_clock),
    .reset(stealServers_30_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_30_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_30_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_30_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_30_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_30_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_30_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_30_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_30_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_30_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_30_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_30_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_30_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_30_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_30_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_30_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_30_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_30_io_connQ_pop_bits)
  );
  stealServer stealServers_31 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_31_clock),
    .reset(stealServers_31_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_31_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_31_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_31_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_31_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_31_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_31_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_31_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_31_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_31_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_31_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_31_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_31_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_31_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_31_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_31_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_31_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_31_io_connQ_pop_bits)
  );
  stealServer stealServers_32 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_32_clock),
    .reset(stealServers_32_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_32_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_32_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_32_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_32_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_32_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_32_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_32_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_32_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_32_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_32_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_32_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_32_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_32_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_32_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_32_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_32_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_32_io_connQ_pop_bits)
  );
  stealServer stealServers_33 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_33_clock),
    .reset(stealServers_33_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_33_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_33_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_33_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_33_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_33_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_33_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_33_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_33_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_33_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_33_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_33_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_33_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_33_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_33_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_33_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_33_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_33_io_connQ_pop_bits)
  );
  stealServer stealServers_34 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_34_clock),
    .reset(stealServers_34_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_34_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_34_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_34_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_34_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_34_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_34_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_34_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_34_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_34_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_34_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_34_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_34_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_34_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_34_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_34_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_34_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_34_io_connQ_pop_bits)
  );
  stealServer stealServers_35 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_35_clock),
    .reset(stealServers_35_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_35_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_35_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_35_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_35_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_35_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_35_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_35_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_35_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_35_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_35_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_35_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_35_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_35_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_35_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_35_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_35_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_35_io_connQ_pop_bits)
  );
  stealServer stealServers_36 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_36_clock),
    .reset(stealServers_36_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_36_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_36_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_36_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_36_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_36_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_36_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_36_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_36_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_36_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_36_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_36_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_36_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_36_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_36_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_36_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_36_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_36_io_connQ_pop_bits)
  );
  stealServer stealServers_37 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_37_clock),
    .reset(stealServers_37_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_37_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_37_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_37_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_37_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_37_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_37_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_37_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_37_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_37_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_37_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_37_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_37_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_37_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_37_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_37_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_37_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_37_io_connQ_pop_bits)
  );
  stealServer stealServers_38 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_38_clock),
    .reset(stealServers_38_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_38_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_38_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_38_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_38_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_38_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_38_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_38_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_38_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_38_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_38_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_38_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_38_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_38_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_38_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_38_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_38_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_38_io_connQ_pop_bits)
  );
  stealServer stealServers_39 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_39_clock),
    .reset(stealServers_39_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_39_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_39_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_39_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_39_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_39_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_39_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_39_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_39_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_39_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_39_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_39_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_39_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_39_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_39_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_39_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_39_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_39_io_connQ_pop_bits)
  );
  stealServer stealServers_40 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_40_clock),
    .reset(stealServers_40_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_40_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_40_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_40_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_40_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_40_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_40_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_40_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_40_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_40_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_40_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_40_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_40_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_40_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_40_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_40_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_40_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_40_io_connQ_pop_bits)
  );
  stealServer stealServers_41 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_41_clock),
    .reset(stealServers_41_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_41_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_41_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_41_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_41_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_41_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_41_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_41_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_41_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_41_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_41_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_41_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_41_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_41_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_41_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_41_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_41_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_41_io_connQ_pop_bits)
  );
  stealServer stealServers_42 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_42_clock),
    .reset(stealServers_42_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_42_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_42_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_42_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_42_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_42_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_42_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_42_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_42_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_42_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_42_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_42_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_42_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_42_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_42_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_42_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_42_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_42_io_connQ_pop_bits)
  );
  stealServer stealServers_43 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_43_clock),
    .reset(stealServers_43_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_43_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_43_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_43_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_43_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_43_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_43_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_43_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_43_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_43_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_43_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_43_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_43_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_43_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_43_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_43_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_43_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_43_io_connQ_pop_bits)
  );
  stealServer stealServers_44 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_44_clock),
    .reset(stealServers_44_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_44_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_44_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_44_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_44_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_44_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_44_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_44_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_44_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_44_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_44_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_44_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_44_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_44_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_44_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_44_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_44_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_44_io_connQ_pop_bits)
  );
  stealServer stealServers_45 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_45_clock),
    .reset(stealServers_45_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_45_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_45_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_45_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_45_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_45_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_45_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_45_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_45_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_45_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_45_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_45_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_45_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_45_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_45_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_45_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_45_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_45_io_connQ_pop_bits)
  );
  stealServer stealServers_46 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_46_clock),
    .reset(stealServers_46_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_46_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_46_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_46_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_46_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_46_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_46_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_46_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_46_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_46_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_46_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_46_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_46_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_46_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_46_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_46_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_46_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_46_io_connQ_pop_bits)
  );
  stealServer stealServers_47 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_47_clock),
    .reset(stealServers_47_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_47_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_47_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_47_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_47_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_47_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_47_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_47_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_47_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_47_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_47_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_47_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_47_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_47_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_47_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_47_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_47_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_47_io_connQ_pop_bits)
  );
  stealServer stealServers_48 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_48_clock),
    .reset(stealServers_48_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_48_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_48_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_48_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_48_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_48_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_48_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_48_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_48_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_48_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_48_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_48_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_48_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_48_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_48_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_48_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_48_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_48_io_connQ_pop_bits)
  );
  stealServer stealServers_49 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_49_clock),
    .reset(stealServers_49_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_49_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_49_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_49_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_49_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_49_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_49_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_49_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_49_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_49_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_49_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_49_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_49_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_49_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_49_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_49_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_49_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_49_io_connQ_pop_bits)
  );
  stealServer stealServers_50 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_50_clock),
    .reset(stealServers_50_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_50_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_50_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_50_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_50_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_50_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_50_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_50_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_50_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_50_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_50_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_50_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_50_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_50_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_50_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_50_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_50_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_50_io_connQ_pop_bits)
  );
  stealServer stealServers_51 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_51_clock),
    .reset(stealServers_51_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_51_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_51_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_51_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_51_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_51_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_51_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_51_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_51_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_51_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_51_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_51_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_51_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_51_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_51_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_51_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_51_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_51_io_connQ_pop_bits)
  );
  stealServer stealServers_52 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_52_clock),
    .reset(stealServers_52_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_52_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_52_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_52_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_52_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_52_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_52_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_52_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_52_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_52_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_52_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_52_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_52_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_52_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_52_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_52_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_52_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_52_io_connQ_pop_bits)
  );
  stealServer stealServers_53 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_53_clock),
    .reset(stealServers_53_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_53_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_53_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_53_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_53_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_53_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_53_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_53_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_53_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_53_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_53_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_53_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_53_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_53_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_53_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_53_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_53_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_53_io_connQ_pop_bits)
  );
  stealServer stealServers_54 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_54_clock),
    .reset(stealServers_54_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_54_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_54_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_54_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_54_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_54_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_54_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_54_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_54_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_54_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_54_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_54_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_54_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_54_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_54_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_54_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_54_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_54_io_connQ_pop_bits)
  );
  stealServer stealServers_55 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_55_clock),
    .reset(stealServers_55_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_55_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_55_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_55_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_55_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_55_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_55_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_55_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_55_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_55_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_55_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_55_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_55_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_55_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_55_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_55_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_55_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_55_io_connQ_pop_bits)
  );
  stealServer stealServers_56 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_56_clock),
    .reset(stealServers_56_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_56_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_56_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_56_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_56_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_56_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_56_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_56_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_56_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_56_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_56_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_56_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_56_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_56_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_56_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_56_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_56_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_56_io_connQ_pop_bits)
  );
  stealServer stealServers_57 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_57_clock),
    .reset(stealServers_57_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_57_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_57_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_57_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_57_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_57_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_57_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_57_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_57_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_57_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_57_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_57_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_57_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_57_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_57_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_57_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_57_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_57_io_connQ_pop_bits)
  );
  stealServer stealServers_58 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_58_clock),
    .reset(stealServers_58_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_58_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_58_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_58_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_58_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_58_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_58_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_58_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_58_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_58_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_58_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_58_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_58_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_58_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_58_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_58_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_58_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_58_io_connQ_pop_bits)
  );
  stealServer stealServers_59 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_59_clock),
    .reset(stealServers_59_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_59_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_59_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_59_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_59_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_59_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_59_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_59_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_59_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_59_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_59_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_59_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_59_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_59_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_59_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_59_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_59_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_59_io_connQ_pop_bits)
  );
  stealServer stealServers_60 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_60_clock),
    .reset(stealServers_60_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_60_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_60_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_60_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_60_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_60_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_60_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_60_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_60_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_60_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_60_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_60_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_60_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_60_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_60_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_60_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_60_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_60_io_connQ_pop_bits)
  );
  stealServer stealServers_61 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_61_clock),
    .reset(stealServers_61_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_61_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_61_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_61_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_61_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_61_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_61_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_61_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_61_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_61_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_61_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_61_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_61_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_61_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_61_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_61_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_61_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_61_io_connQ_pop_bits)
  );
  stealServer stealServers_62 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_62_clock),
    .reset(stealServers_62_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_62_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_62_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_62_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_62_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_62_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_62_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_62_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_62_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_62_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_62_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_62_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_62_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_62_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_62_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_62_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_62_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_62_io_connQ_pop_bits)
  );
  stealServer stealServers_63 ( // @[stealNW_TQ.scala 54:49]
    .clock(stealServers_63_clock),
    .reset(stealServers_63_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(stealServers_63_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(stealServers_63_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_ctrl_stealReq_ready(stealServers_63_io_connNetwork_ctrl_stealReq_ready),
    .io_connNetwork_ctrl_stealReq_valid(stealServers_63_io_connNetwork_ctrl_stealReq_valid),
    .io_connNetwork_data_availableTask_ready(stealServers_63_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(stealServers_63_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(stealServers_63_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(stealServers_63_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(stealServers_63_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(stealServers_63_io_connNetwork_data_qOutTask_bits),
    .io_connQ_currLength(stealServers_63_io_connQ_currLength),
    .io_connQ_push_ready(stealServers_63_io_connQ_push_ready),
    .io_connQ_push_valid(stealServers_63_io_connQ_push_valid),
    .io_connQ_push_bits(stealServers_63_io_connQ_push_bits),
    .io_connQ_pop_ready(stealServers_63_io_connQ_pop_ready),
    .io_connQ_pop_valid(stealServers_63_io_connQ_pop_valid),
    .io_connQ_pop_bits(stealServers_63_io_connQ_pop_bits)
  );
  hw_deque taskQueues_0 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_0_clock),
    .reset(taskQueues_0_reset),
    .io_connVec_0_push_ready(taskQueues_0_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_0_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_0_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_0_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_0_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_0_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_0_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_0_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_0_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_0_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_0_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_0_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_0_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_1 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_1_clock),
    .reset(taskQueues_1_reset),
    .io_connVec_0_push_ready(taskQueues_1_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_1_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_1_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_1_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_1_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_1_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_1_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_1_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_1_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_1_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_1_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_1_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_1_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_2 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_2_clock),
    .reset(taskQueues_2_reset),
    .io_connVec_0_push_ready(taskQueues_2_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_2_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_2_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_2_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_2_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_2_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_2_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_2_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_2_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_2_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_2_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_2_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_2_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_3 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_3_clock),
    .reset(taskQueues_3_reset),
    .io_connVec_0_push_ready(taskQueues_3_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_3_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_3_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_3_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_3_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_3_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_3_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_3_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_3_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_3_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_3_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_3_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_3_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_4 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_4_clock),
    .reset(taskQueues_4_reset),
    .io_connVec_0_push_ready(taskQueues_4_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_4_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_4_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_4_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_4_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_4_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_4_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_4_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_4_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_4_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_4_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_4_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_4_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_5 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_5_clock),
    .reset(taskQueues_5_reset),
    .io_connVec_0_push_ready(taskQueues_5_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_5_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_5_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_5_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_5_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_5_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_5_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_5_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_5_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_5_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_5_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_5_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_5_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_6 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_6_clock),
    .reset(taskQueues_6_reset),
    .io_connVec_0_push_ready(taskQueues_6_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_6_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_6_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_6_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_6_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_6_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_6_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_6_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_6_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_6_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_6_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_6_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_6_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_7 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_7_clock),
    .reset(taskQueues_7_reset),
    .io_connVec_0_push_ready(taskQueues_7_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_7_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_7_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_7_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_7_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_7_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_7_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_7_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_7_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_7_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_7_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_7_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_7_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_8 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_8_clock),
    .reset(taskQueues_8_reset),
    .io_connVec_0_push_ready(taskQueues_8_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_8_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_8_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_8_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_8_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_8_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_8_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_8_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_8_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_8_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_8_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_8_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_8_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_9 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_9_clock),
    .reset(taskQueues_9_reset),
    .io_connVec_0_push_ready(taskQueues_9_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_9_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_9_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_9_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_9_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_9_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_9_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_9_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_9_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_9_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_9_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_9_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_9_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_10 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_10_clock),
    .reset(taskQueues_10_reset),
    .io_connVec_0_push_ready(taskQueues_10_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_10_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_10_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_10_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_10_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_10_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_10_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_10_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_10_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_10_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_10_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_10_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_10_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_11 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_11_clock),
    .reset(taskQueues_11_reset),
    .io_connVec_0_push_ready(taskQueues_11_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_11_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_11_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_11_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_11_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_11_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_11_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_11_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_11_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_11_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_11_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_11_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_11_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_12 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_12_clock),
    .reset(taskQueues_12_reset),
    .io_connVec_0_push_ready(taskQueues_12_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_12_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_12_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_12_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_12_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_12_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_12_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_12_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_12_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_12_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_12_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_12_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_12_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_13 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_13_clock),
    .reset(taskQueues_13_reset),
    .io_connVec_0_push_ready(taskQueues_13_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_13_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_13_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_13_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_13_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_13_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_13_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_13_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_13_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_13_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_13_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_13_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_13_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_14 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_14_clock),
    .reset(taskQueues_14_reset),
    .io_connVec_0_push_ready(taskQueues_14_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_14_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_14_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_14_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_14_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_14_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_14_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_14_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_14_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_14_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_14_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_14_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_14_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_15 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_15_clock),
    .reset(taskQueues_15_reset),
    .io_connVec_0_push_ready(taskQueues_15_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_15_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_15_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_15_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_15_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_15_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_15_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_15_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_15_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_15_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_15_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_15_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_15_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_16 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_16_clock),
    .reset(taskQueues_16_reset),
    .io_connVec_0_push_ready(taskQueues_16_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_16_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_16_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_16_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_16_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_16_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_16_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_16_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_16_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_16_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_16_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_16_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_16_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_17 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_17_clock),
    .reset(taskQueues_17_reset),
    .io_connVec_0_push_ready(taskQueues_17_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_17_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_17_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_17_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_17_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_17_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_17_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_17_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_17_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_17_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_17_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_17_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_17_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_18 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_18_clock),
    .reset(taskQueues_18_reset),
    .io_connVec_0_push_ready(taskQueues_18_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_18_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_18_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_18_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_18_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_18_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_18_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_18_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_18_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_18_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_18_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_18_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_18_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_19 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_19_clock),
    .reset(taskQueues_19_reset),
    .io_connVec_0_push_ready(taskQueues_19_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_19_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_19_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_19_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_19_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_19_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_19_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_19_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_19_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_19_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_19_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_19_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_19_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_20 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_20_clock),
    .reset(taskQueues_20_reset),
    .io_connVec_0_push_ready(taskQueues_20_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_20_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_20_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_20_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_20_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_20_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_20_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_20_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_20_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_20_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_20_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_20_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_20_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_21 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_21_clock),
    .reset(taskQueues_21_reset),
    .io_connVec_0_push_ready(taskQueues_21_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_21_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_21_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_21_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_21_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_21_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_21_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_21_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_21_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_21_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_21_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_21_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_21_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_22 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_22_clock),
    .reset(taskQueues_22_reset),
    .io_connVec_0_push_ready(taskQueues_22_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_22_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_22_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_22_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_22_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_22_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_22_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_22_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_22_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_22_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_22_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_22_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_22_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_23 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_23_clock),
    .reset(taskQueues_23_reset),
    .io_connVec_0_push_ready(taskQueues_23_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_23_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_23_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_23_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_23_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_23_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_23_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_23_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_23_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_23_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_23_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_23_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_23_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_24 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_24_clock),
    .reset(taskQueues_24_reset),
    .io_connVec_0_push_ready(taskQueues_24_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_24_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_24_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_24_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_24_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_24_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_24_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_24_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_24_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_24_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_24_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_24_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_24_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_25 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_25_clock),
    .reset(taskQueues_25_reset),
    .io_connVec_0_push_ready(taskQueues_25_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_25_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_25_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_25_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_25_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_25_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_25_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_25_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_25_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_25_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_25_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_25_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_25_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_26 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_26_clock),
    .reset(taskQueues_26_reset),
    .io_connVec_0_push_ready(taskQueues_26_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_26_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_26_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_26_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_26_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_26_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_26_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_26_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_26_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_26_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_26_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_26_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_26_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_27 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_27_clock),
    .reset(taskQueues_27_reset),
    .io_connVec_0_push_ready(taskQueues_27_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_27_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_27_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_27_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_27_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_27_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_27_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_27_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_27_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_27_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_27_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_27_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_27_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_28 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_28_clock),
    .reset(taskQueues_28_reset),
    .io_connVec_0_push_ready(taskQueues_28_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_28_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_28_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_28_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_28_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_28_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_28_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_28_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_28_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_28_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_28_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_28_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_28_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_29 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_29_clock),
    .reset(taskQueues_29_reset),
    .io_connVec_0_push_ready(taskQueues_29_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_29_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_29_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_29_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_29_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_29_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_29_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_29_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_29_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_29_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_29_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_29_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_29_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_30 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_30_clock),
    .reset(taskQueues_30_reset),
    .io_connVec_0_push_ready(taskQueues_30_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_30_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_30_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_30_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_30_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_30_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_30_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_30_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_30_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_30_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_30_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_30_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_30_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_31 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_31_clock),
    .reset(taskQueues_31_reset),
    .io_connVec_0_push_ready(taskQueues_31_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_31_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_31_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_31_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_31_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_31_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_31_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_31_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_31_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_31_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_31_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_31_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_31_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_32 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_32_clock),
    .reset(taskQueues_32_reset),
    .io_connVec_0_push_ready(taskQueues_32_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_32_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_32_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_32_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_32_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_32_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_32_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_32_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_32_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_32_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_32_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_32_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_32_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_33 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_33_clock),
    .reset(taskQueues_33_reset),
    .io_connVec_0_push_ready(taskQueues_33_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_33_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_33_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_33_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_33_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_33_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_33_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_33_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_33_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_33_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_33_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_33_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_33_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_34 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_34_clock),
    .reset(taskQueues_34_reset),
    .io_connVec_0_push_ready(taskQueues_34_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_34_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_34_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_34_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_34_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_34_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_34_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_34_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_34_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_34_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_34_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_34_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_34_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_35 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_35_clock),
    .reset(taskQueues_35_reset),
    .io_connVec_0_push_ready(taskQueues_35_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_35_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_35_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_35_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_35_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_35_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_35_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_35_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_35_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_35_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_35_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_35_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_35_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_36 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_36_clock),
    .reset(taskQueues_36_reset),
    .io_connVec_0_push_ready(taskQueues_36_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_36_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_36_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_36_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_36_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_36_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_36_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_36_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_36_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_36_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_36_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_36_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_36_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_37 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_37_clock),
    .reset(taskQueues_37_reset),
    .io_connVec_0_push_ready(taskQueues_37_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_37_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_37_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_37_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_37_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_37_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_37_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_37_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_37_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_37_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_37_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_37_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_37_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_38 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_38_clock),
    .reset(taskQueues_38_reset),
    .io_connVec_0_push_ready(taskQueues_38_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_38_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_38_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_38_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_38_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_38_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_38_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_38_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_38_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_38_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_38_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_38_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_38_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_39 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_39_clock),
    .reset(taskQueues_39_reset),
    .io_connVec_0_push_ready(taskQueues_39_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_39_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_39_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_39_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_39_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_39_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_39_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_39_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_39_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_39_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_39_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_39_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_39_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_40 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_40_clock),
    .reset(taskQueues_40_reset),
    .io_connVec_0_push_ready(taskQueues_40_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_40_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_40_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_40_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_40_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_40_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_40_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_40_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_40_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_40_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_40_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_40_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_40_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_41 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_41_clock),
    .reset(taskQueues_41_reset),
    .io_connVec_0_push_ready(taskQueues_41_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_41_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_41_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_41_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_41_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_41_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_41_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_41_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_41_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_41_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_41_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_41_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_41_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_42 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_42_clock),
    .reset(taskQueues_42_reset),
    .io_connVec_0_push_ready(taskQueues_42_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_42_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_42_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_42_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_42_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_42_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_42_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_42_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_42_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_42_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_42_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_42_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_42_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_43 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_43_clock),
    .reset(taskQueues_43_reset),
    .io_connVec_0_push_ready(taskQueues_43_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_43_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_43_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_43_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_43_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_43_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_43_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_43_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_43_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_43_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_43_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_43_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_43_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_44 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_44_clock),
    .reset(taskQueues_44_reset),
    .io_connVec_0_push_ready(taskQueues_44_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_44_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_44_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_44_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_44_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_44_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_44_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_44_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_44_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_44_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_44_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_44_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_44_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_45 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_45_clock),
    .reset(taskQueues_45_reset),
    .io_connVec_0_push_ready(taskQueues_45_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_45_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_45_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_45_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_45_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_45_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_45_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_45_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_45_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_45_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_45_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_45_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_45_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_46 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_46_clock),
    .reset(taskQueues_46_reset),
    .io_connVec_0_push_ready(taskQueues_46_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_46_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_46_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_46_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_46_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_46_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_46_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_46_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_46_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_46_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_46_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_46_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_46_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_47 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_47_clock),
    .reset(taskQueues_47_reset),
    .io_connVec_0_push_ready(taskQueues_47_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_47_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_47_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_47_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_47_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_47_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_47_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_47_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_47_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_47_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_47_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_47_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_47_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_48 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_48_clock),
    .reset(taskQueues_48_reset),
    .io_connVec_0_push_ready(taskQueues_48_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_48_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_48_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_48_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_48_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_48_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_48_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_48_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_48_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_48_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_48_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_48_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_48_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_49 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_49_clock),
    .reset(taskQueues_49_reset),
    .io_connVec_0_push_ready(taskQueues_49_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_49_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_49_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_49_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_49_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_49_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_49_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_49_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_49_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_49_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_49_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_49_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_49_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_50 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_50_clock),
    .reset(taskQueues_50_reset),
    .io_connVec_0_push_ready(taskQueues_50_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_50_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_50_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_50_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_50_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_50_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_50_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_50_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_50_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_50_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_50_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_50_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_50_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_51 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_51_clock),
    .reset(taskQueues_51_reset),
    .io_connVec_0_push_ready(taskQueues_51_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_51_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_51_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_51_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_51_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_51_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_51_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_51_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_51_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_51_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_51_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_51_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_51_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_52 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_52_clock),
    .reset(taskQueues_52_reset),
    .io_connVec_0_push_ready(taskQueues_52_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_52_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_52_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_52_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_52_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_52_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_52_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_52_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_52_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_52_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_52_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_52_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_52_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_53 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_53_clock),
    .reset(taskQueues_53_reset),
    .io_connVec_0_push_ready(taskQueues_53_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_53_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_53_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_53_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_53_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_53_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_53_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_53_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_53_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_53_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_53_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_53_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_53_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_54 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_54_clock),
    .reset(taskQueues_54_reset),
    .io_connVec_0_push_ready(taskQueues_54_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_54_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_54_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_54_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_54_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_54_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_54_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_54_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_54_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_54_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_54_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_54_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_54_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_55 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_55_clock),
    .reset(taskQueues_55_reset),
    .io_connVec_0_push_ready(taskQueues_55_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_55_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_55_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_55_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_55_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_55_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_55_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_55_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_55_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_55_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_55_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_55_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_55_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_56 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_56_clock),
    .reset(taskQueues_56_reset),
    .io_connVec_0_push_ready(taskQueues_56_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_56_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_56_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_56_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_56_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_56_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_56_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_56_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_56_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_56_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_56_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_56_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_56_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_57 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_57_clock),
    .reset(taskQueues_57_reset),
    .io_connVec_0_push_ready(taskQueues_57_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_57_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_57_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_57_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_57_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_57_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_57_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_57_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_57_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_57_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_57_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_57_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_57_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_58 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_58_clock),
    .reset(taskQueues_58_reset),
    .io_connVec_0_push_ready(taskQueues_58_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_58_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_58_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_58_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_58_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_58_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_58_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_58_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_58_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_58_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_58_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_58_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_58_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_59 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_59_clock),
    .reset(taskQueues_59_reset),
    .io_connVec_0_push_ready(taskQueues_59_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_59_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_59_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_59_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_59_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_59_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_59_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_59_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_59_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_59_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_59_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_59_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_59_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_60 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_60_clock),
    .reset(taskQueues_60_reset),
    .io_connVec_0_push_ready(taskQueues_60_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_60_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_60_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_60_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_60_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_60_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_60_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_60_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_60_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_60_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_60_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_60_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_60_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_61 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_61_clock),
    .reset(taskQueues_61_reset),
    .io_connVec_0_push_ready(taskQueues_61_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_61_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_61_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_61_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_61_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_61_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_61_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_61_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_61_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_61_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_61_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_61_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_61_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_62 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_62_clock),
    .reset(taskQueues_62_reset),
    .io_connVec_0_push_ready(taskQueues_62_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_62_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_62_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_62_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_62_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_62_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_62_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_62_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_62_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_62_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_62_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_62_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_62_io_connVec_1_pop_bits)
  );
  hw_deque taskQueues_63 ( // @[stealNW_TQ.scala 58:49]
    .clock(taskQueues_63_clock),
    .reset(taskQueues_63_reset),
    .io_connVec_0_push_ready(taskQueues_63_io_connVec_0_push_ready),
    .io_connVec_0_push_valid(taskQueues_63_io_connVec_0_push_valid),
    .io_connVec_0_push_bits(taskQueues_63_io_connVec_0_push_bits),
    .io_connVec_0_pop_ready(taskQueues_63_io_connVec_0_pop_ready),
    .io_connVec_0_pop_valid(taskQueues_63_io_connVec_0_pop_valid),
    .io_connVec_0_pop_bits(taskQueues_63_io_connVec_0_pop_bits),
    .io_connVec_1_currLength(taskQueues_63_io_connVec_1_currLength),
    .io_connVec_1_push_ready(taskQueues_63_io_connVec_1_push_ready),
    .io_connVec_1_push_valid(taskQueues_63_io_connVec_1_push_valid),
    .io_connVec_1_push_bits(taskQueues_63_io_connVec_1_push_bits),
    .io_connVec_1_pop_ready(taskQueues_63_io_connVec_1_pop_ready),
    .io_connVec_1_pop_valid(taskQueues_63_io_connVec_1_pop_valid),
    .io_connVec_1_pop_bits(taskQueues_63_io_connVec_1_pop_bits)
  );
  assign io_connPE_0_push_ready = taskQueues_0_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_0_pop_valid = taskQueues_0_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_0_pop_bits = taskQueues_0_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_1_push_ready = taskQueues_1_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_1_pop_valid = taskQueues_1_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_1_pop_bits = taskQueues_1_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_2_push_ready = taskQueues_2_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_2_pop_valid = taskQueues_2_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_2_pop_bits = taskQueues_2_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_3_push_ready = taskQueues_3_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_3_pop_valid = taskQueues_3_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_3_pop_bits = taskQueues_3_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_4_push_ready = taskQueues_4_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_4_pop_valid = taskQueues_4_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_4_pop_bits = taskQueues_4_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_5_push_ready = taskQueues_5_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_5_pop_valid = taskQueues_5_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_5_pop_bits = taskQueues_5_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_6_push_ready = taskQueues_6_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_6_pop_valid = taskQueues_6_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_6_pop_bits = taskQueues_6_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_7_push_ready = taskQueues_7_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_7_pop_valid = taskQueues_7_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_7_pop_bits = taskQueues_7_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_8_push_ready = taskQueues_8_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_8_pop_valid = taskQueues_8_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_8_pop_bits = taskQueues_8_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_9_push_ready = taskQueues_9_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_9_pop_valid = taskQueues_9_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_9_pop_bits = taskQueues_9_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_10_push_ready = taskQueues_10_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_10_pop_valid = taskQueues_10_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_10_pop_bits = taskQueues_10_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_11_push_ready = taskQueues_11_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_11_pop_valid = taskQueues_11_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_11_pop_bits = taskQueues_11_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_12_push_ready = taskQueues_12_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_12_pop_valid = taskQueues_12_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_12_pop_bits = taskQueues_12_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_13_push_ready = taskQueues_13_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_13_pop_valid = taskQueues_13_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_13_pop_bits = taskQueues_13_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_14_push_ready = taskQueues_14_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_14_pop_valid = taskQueues_14_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_14_pop_bits = taskQueues_14_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_15_push_ready = taskQueues_15_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_15_pop_valid = taskQueues_15_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_15_pop_bits = taskQueues_15_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_16_push_ready = taskQueues_16_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_16_pop_valid = taskQueues_16_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_16_pop_bits = taskQueues_16_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_17_push_ready = taskQueues_17_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_17_pop_valid = taskQueues_17_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_17_pop_bits = taskQueues_17_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_18_push_ready = taskQueues_18_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_18_pop_valid = taskQueues_18_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_18_pop_bits = taskQueues_18_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_19_push_ready = taskQueues_19_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_19_pop_valid = taskQueues_19_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_19_pop_bits = taskQueues_19_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_20_push_ready = taskQueues_20_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_20_pop_valid = taskQueues_20_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_20_pop_bits = taskQueues_20_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_21_push_ready = taskQueues_21_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_21_pop_valid = taskQueues_21_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_21_pop_bits = taskQueues_21_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_22_push_ready = taskQueues_22_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_22_pop_valid = taskQueues_22_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_22_pop_bits = taskQueues_22_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_23_push_ready = taskQueues_23_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_23_pop_valid = taskQueues_23_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_23_pop_bits = taskQueues_23_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_24_push_ready = taskQueues_24_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_24_pop_valid = taskQueues_24_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_24_pop_bits = taskQueues_24_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_25_push_ready = taskQueues_25_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_25_pop_valid = taskQueues_25_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_25_pop_bits = taskQueues_25_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_26_push_ready = taskQueues_26_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_26_pop_valid = taskQueues_26_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_26_pop_bits = taskQueues_26_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_27_push_ready = taskQueues_27_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_27_pop_valid = taskQueues_27_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_27_pop_bits = taskQueues_27_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_28_push_ready = taskQueues_28_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_28_pop_valid = taskQueues_28_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_28_pop_bits = taskQueues_28_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_29_push_ready = taskQueues_29_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_29_pop_valid = taskQueues_29_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_29_pop_bits = taskQueues_29_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_30_push_ready = taskQueues_30_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_30_pop_valid = taskQueues_30_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_30_pop_bits = taskQueues_30_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_31_push_ready = taskQueues_31_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_31_pop_valid = taskQueues_31_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_31_pop_bits = taskQueues_31_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_32_push_ready = taskQueues_32_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_32_pop_valid = taskQueues_32_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_32_pop_bits = taskQueues_32_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_33_push_ready = taskQueues_33_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_33_pop_valid = taskQueues_33_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_33_pop_bits = taskQueues_33_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_34_push_ready = taskQueues_34_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_34_pop_valid = taskQueues_34_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_34_pop_bits = taskQueues_34_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_35_push_ready = taskQueues_35_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_35_pop_valid = taskQueues_35_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_35_pop_bits = taskQueues_35_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_36_push_ready = taskQueues_36_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_36_pop_valid = taskQueues_36_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_36_pop_bits = taskQueues_36_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_37_push_ready = taskQueues_37_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_37_pop_valid = taskQueues_37_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_37_pop_bits = taskQueues_37_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_38_push_ready = taskQueues_38_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_38_pop_valid = taskQueues_38_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_38_pop_bits = taskQueues_38_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_39_push_ready = taskQueues_39_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_39_pop_valid = taskQueues_39_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_39_pop_bits = taskQueues_39_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_40_push_ready = taskQueues_40_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_40_pop_valid = taskQueues_40_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_40_pop_bits = taskQueues_40_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_41_push_ready = taskQueues_41_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_41_pop_valid = taskQueues_41_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_41_pop_bits = taskQueues_41_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_42_push_ready = taskQueues_42_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_42_pop_valid = taskQueues_42_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_42_pop_bits = taskQueues_42_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_43_push_ready = taskQueues_43_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_43_pop_valid = taskQueues_43_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_43_pop_bits = taskQueues_43_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_44_push_ready = taskQueues_44_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_44_pop_valid = taskQueues_44_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_44_pop_bits = taskQueues_44_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_45_push_ready = taskQueues_45_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_45_pop_valid = taskQueues_45_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_45_pop_bits = taskQueues_45_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_46_push_ready = taskQueues_46_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_46_pop_valid = taskQueues_46_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_46_pop_bits = taskQueues_46_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_47_push_ready = taskQueues_47_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_47_pop_valid = taskQueues_47_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_47_pop_bits = taskQueues_47_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_48_push_ready = taskQueues_48_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_48_pop_valid = taskQueues_48_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_48_pop_bits = taskQueues_48_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_49_push_ready = taskQueues_49_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_49_pop_valid = taskQueues_49_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_49_pop_bits = taskQueues_49_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_50_push_ready = taskQueues_50_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_50_pop_valid = taskQueues_50_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_50_pop_bits = taskQueues_50_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_51_push_ready = taskQueues_51_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_51_pop_valid = taskQueues_51_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_51_pop_bits = taskQueues_51_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_52_push_ready = taskQueues_52_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_52_pop_valid = taskQueues_52_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_52_pop_bits = taskQueues_52_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_53_push_ready = taskQueues_53_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_53_pop_valid = taskQueues_53_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_53_pop_bits = taskQueues_53_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_54_push_ready = taskQueues_54_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_54_pop_valid = taskQueues_54_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_54_pop_bits = taskQueues_54_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_55_push_ready = taskQueues_55_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_55_pop_valid = taskQueues_55_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_55_pop_bits = taskQueues_55_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_56_push_ready = taskQueues_56_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_56_pop_valid = taskQueues_56_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_56_pop_bits = taskQueues_56_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_57_push_ready = taskQueues_57_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_57_pop_valid = taskQueues_57_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_57_pop_bits = taskQueues_57_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_58_push_ready = taskQueues_58_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_58_pop_valid = taskQueues_58_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_58_pop_bits = taskQueues_58_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_59_push_ready = taskQueues_59_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_59_pop_valid = taskQueues_59_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_59_pop_bits = taskQueues_59_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_60_push_ready = taskQueues_60_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_60_pop_valid = taskQueues_60_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_60_pop_bits = taskQueues_60_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_61_push_ready = taskQueues_61_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_61_pop_valid = taskQueues_61_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_61_pop_bits = taskQueues_61_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_62_push_ready = taskQueues_62_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_62_pop_valid = taskQueues_62_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_62_pop_bits = taskQueues_62_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_63_push_ready = taskQueues_63_io_connVec_0_push_ready; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_63_pop_valid = taskQueues_63_io_connVec_0_pop_valid; // @[stealNW_TQ.scala 62:37]
  assign io_connPE_63_pop_bits = taskQueues_63_io_connVec_0_pop_bits; // @[stealNW_TQ.scala 62:37]
  assign io_connVSS_0_ctrl_serveStealReq_ready = stealNet_io_connSS_2_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 107:44]
  assign io_connVSS_0_data_availableTask_valid = stealNet_io_connSS_0_data_availableTask_valid; // @[stealNW_TQ.scala 87:44]
  assign io_connVSS_0_data_availableTask_bits = stealNet_io_connSS_0_data_availableTask_bits; // @[stealNW_TQ.scala 87:44]
  assign io_connVSS_0_data_qOutTask_ready = stealNet_io_connSS_0_data_qOutTask_ready; // @[stealNW_TQ.scala 87:44]
  assign io_connVAS_0_ctrl_serveStealReq_ready = stealNet_io_connSS_0_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 104:44]
  assign io_connVAS_0_data_qOutTask_ready = stealNet_io_connSS_1_data_qOutTask_ready; // @[stealNW_TQ.scala 90:44]
  assign io_connVAS_1_ctrl_serveStealReq_ready = stealNet_io_connSS_1_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 104:44]
  assign io_connVAS_1_data_qOutTask_ready = stealNet_io_connSS_2_data_qOutTask_ready; // @[stealNW_TQ.scala 90:44]
  assign io_ntwDataUnitOccupancyVSS_0 = stealNet_io_ntwDataUnitOccupancyVSS_0; // @[stealNW_TQ.scala 145:48]
  assign stealNet_clock = clock;
  assign stealNet_reset = reset;
  assign stealNet_io_connSS_0_ctrl_serveStealReq_valid = io_connVAS_0_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 104:44]
  assign stealNet_io_connSS_0_data_availableTask_ready = io_connVSS_0_data_availableTask_ready; // @[stealNW_TQ.scala 87:44]
  assign stealNet_io_connSS_0_data_qOutTask_valid = io_connVSS_0_data_qOutTask_valid; // @[stealNW_TQ.scala 87:44]
  assign stealNet_io_connSS_0_data_qOutTask_bits = io_connVSS_0_data_qOutTask_bits; // @[stealNW_TQ.scala 87:44]
  assign stealNet_io_connSS_1_ctrl_serveStealReq_valid = io_connVAS_1_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 104:44]
  assign stealNet_io_connSS_1_data_qOutTask_valid = io_connVAS_0_data_qOutTask_valid; // @[stealNW_TQ.scala 90:44]
  assign stealNet_io_connSS_1_data_qOutTask_bits = io_connVAS_0_data_qOutTask_bits; // @[stealNW_TQ.scala 90:44]
  assign stealNet_io_connSS_2_ctrl_serveStealReq_valid = io_connVSS_0_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 107:44]
  assign stealNet_io_connSS_2_data_qOutTask_valid = io_connVAS_1_data_qOutTask_valid; // @[stealNW_TQ.scala 90:44]
  assign stealNet_io_connSS_2_data_qOutTask_bits = io_connVAS_1_data_qOutTask_bits; // @[stealNW_TQ.scala 90:44]
  assign stealNet_io_connSS_3_ctrl_serveStealReq_valid = stealServers_0_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_3_ctrl_stealReq_valid = stealServers_0_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_3_data_availableTask_ready = stealServers_0_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_3_data_qOutTask_valid = stealServers_0_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_3_data_qOutTask_bits = stealServers_0_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_4_ctrl_serveStealReq_valid = stealServers_1_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_4_ctrl_stealReq_valid = stealServers_1_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_4_data_availableTask_ready = stealServers_1_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_4_data_qOutTask_valid = stealServers_1_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_4_data_qOutTask_bits = stealServers_1_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_5_ctrl_serveStealReq_valid = stealServers_2_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_5_ctrl_stealReq_valid = stealServers_2_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_5_data_availableTask_ready = stealServers_2_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_5_data_qOutTask_valid = stealServers_2_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_5_data_qOutTask_bits = stealServers_2_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_6_ctrl_serveStealReq_valid = stealServers_3_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_6_ctrl_stealReq_valid = stealServers_3_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_6_data_availableTask_ready = stealServers_3_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_6_data_qOutTask_valid = stealServers_3_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_6_data_qOutTask_bits = stealServers_3_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_7_ctrl_serveStealReq_valid = stealServers_4_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_7_ctrl_stealReq_valid = stealServers_4_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_7_data_availableTask_ready = stealServers_4_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_7_data_qOutTask_valid = stealServers_4_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_7_data_qOutTask_bits = stealServers_4_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_8_ctrl_serveStealReq_valid = stealServers_5_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_8_ctrl_stealReq_valid = stealServers_5_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_8_data_availableTask_ready = stealServers_5_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_8_data_qOutTask_valid = stealServers_5_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_8_data_qOutTask_bits = stealServers_5_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_9_ctrl_serveStealReq_valid = stealServers_6_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_9_ctrl_stealReq_valid = stealServers_6_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_9_data_availableTask_ready = stealServers_6_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_9_data_qOutTask_valid = stealServers_6_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_9_data_qOutTask_bits = stealServers_6_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_10_ctrl_serveStealReq_valid = stealServers_7_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_10_ctrl_stealReq_valid = stealServers_7_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_10_data_availableTask_ready = stealServers_7_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_10_data_qOutTask_valid = stealServers_7_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_10_data_qOutTask_bits = stealServers_7_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_11_ctrl_serveStealReq_valid = stealServers_8_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_11_ctrl_stealReq_valid = stealServers_8_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_11_data_availableTask_ready = stealServers_8_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_11_data_qOutTask_valid = stealServers_8_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_11_data_qOutTask_bits = stealServers_8_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_12_ctrl_serveStealReq_valid = stealServers_9_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_12_ctrl_stealReq_valid = stealServers_9_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_12_data_availableTask_ready = stealServers_9_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_12_data_qOutTask_valid = stealServers_9_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_12_data_qOutTask_bits = stealServers_9_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_13_ctrl_serveStealReq_valid = stealServers_10_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_13_ctrl_stealReq_valid = stealServers_10_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_13_data_availableTask_ready = stealServers_10_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_13_data_qOutTask_valid = stealServers_10_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_13_data_qOutTask_bits = stealServers_10_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_14_ctrl_serveStealReq_valid = stealServers_11_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_14_ctrl_stealReq_valid = stealServers_11_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_14_data_availableTask_ready = stealServers_11_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_14_data_qOutTask_valid = stealServers_11_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_14_data_qOutTask_bits = stealServers_11_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_15_ctrl_serveStealReq_valid = stealServers_12_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_15_ctrl_stealReq_valid = stealServers_12_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_15_data_availableTask_ready = stealServers_12_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_15_data_qOutTask_valid = stealServers_12_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_15_data_qOutTask_bits = stealServers_12_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_16_ctrl_serveStealReq_valid = stealServers_13_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_16_ctrl_stealReq_valid = stealServers_13_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_16_data_availableTask_ready = stealServers_13_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_16_data_qOutTask_valid = stealServers_13_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_16_data_qOutTask_bits = stealServers_13_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_17_ctrl_serveStealReq_valid = stealServers_14_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_17_ctrl_stealReq_valid = stealServers_14_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_17_data_availableTask_ready = stealServers_14_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_17_data_qOutTask_valid = stealServers_14_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_17_data_qOutTask_bits = stealServers_14_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_18_ctrl_serveStealReq_valid = stealServers_15_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_18_ctrl_stealReq_valid = stealServers_15_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_18_data_availableTask_ready = stealServers_15_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_18_data_qOutTask_valid = stealServers_15_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_18_data_qOutTask_bits = stealServers_15_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_19_ctrl_serveStealReq_valid = stealServers_16_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_19_ctrl_stealReq_valid = stealServers_16_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_19_data_availableTask_ready = stealServers_16_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_19_data_qOutTask_valid = stealServers_16_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_19_data_qOutTask_bits = stealServers_16_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_20_ctrl_serveStealReq_valid = stealServers_17_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_20_ctrl_stealReq_valid = stealServers_17_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_20_data_availableTask_ready = stealServers_17_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_20_data_qOutTask_valid = stealServers_17_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_20_data_qOutTask_bits = stealServers_17_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_21_ctrl_serveStealReq_valid = stealServers_18_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_21_ctrl_stealReq_valid = stealServers_18_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_21_data_availableTask_ready = stealServers_18_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_21_data_qOutTask_valid = stealServers_18_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_21_data_qOutTask_bits = stealServers_18_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_22_ctrl_serveStealReq_valid = stealServers_19_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_22_ctrl_stealReq_valid = stealServers_19_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_22_data_availableTask_ready = stealServers_19_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_22_data_qOutTask_valid = stealServers_19_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_22_data_qOutTask_bits = stealServers_19_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_23_ctrl_serveStealReq_valid = stealServers_20_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_23_ctrl_stealReq_valid = stealServers_20_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_23_data_availableTask_ready = stealServers_20_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_23_data_qOutTask_valid = stealServers_20_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_23_data_qOutTask_bits = stealServers_20_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_24_ctrl_serveStealReq_valid = stealServers_21_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_24_ctrl_stealReq_valid = stealServers_21_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_24_data_availableTask_ready = stealServers_21_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_24_data_qOutTask_valid = stealServers_21_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_24_data_qOutTask_bits = stealServers_21_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_25_ctrl_serveStealReq_valid = stealServers_22_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_25_ctrl_stealReq_valid = stealServers_22_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_25_data_availableTask_ready = stealServers_22_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_25_data_qOutTask_valid = stealServers_22_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_25_data_qOutTask_bits = stealServers_22_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_26_ctrl_serveStealReq_valid = stealServers_23_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_26_ctrl_stealReq_valid = stealServers_23_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_26_data_availableTask_ready = stealServers_23_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_26_data_qOutTask_valid = stealServers_23_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_26_data_qOutTask_bits = stealServers_23_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_27_ctrl_serveStealReq_valid = stealServers_24_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_27_ctrl_stealReq_valid = stealServers_24_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_27_data_availableTask_ready = stealServers_24_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_27_data_qOutTask_valid = stealServers_24_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_27_data_qOutTask_bits = stealServers_24_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_28_ctrl_serveStealReq_valid = stealServers_25_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_28_ctrl_stealReq_valid = stealServers_25_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_28_data_availableTask_ready = stealServers_25_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_28_data_qOutTask_valid = stealServers_25_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_28_data_qOutTask_bits = stealServers_25_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_29_ctrl_serveStealReq_valid = stealServers_26_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_29_ctrl_stealReq_valid = stealServers_26_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_29_data_availableTask_ready = stealServers_26_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_29_data_qOutTask_valid = stealServers_26_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_29_data_qOutTask_bits = stealServers_26_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_30_ctrl_serveStealReq_valid = stealServers_27_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_30_ctrl_stealReq_valid = stealServers_27_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_30_data_availableTask_ready = stealServers_27_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_30_data_qOutTask_valid = stealServers_27_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_30_data_qOutTask_bits = stealServers_27_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_31_ctrl_serveStealReq_valid = stealServers_28_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_31_ctrl_stealReq_valid = stealServers_28_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_31_data_availableTask_ready = stealServers_28_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_31_data_qOutTask_valid = stealServers_28_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_31_data_qOutTask_bits = stealServers_28_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_32_ctrl_serveStealReq_valid = stealServers_29_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_32_ctrl_stealReq_valid = stealServers_29_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_32_data_availableTask_ready = stealServers_29_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_32_data_qOutTask_valid = stealServers_29_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_32_data_qOutTask_bits = stealServers_29_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_33_ctrl_serveStealReq_valid = stealServers_30_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_33_ctrl_stealReq_valid = stealServers_30_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_33_data_availableTask_ready = stealServers_30_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_33_data_qOutTask_valid = stealServers_30_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_33_data_qOutTask_bits = stealServers_30_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_34_ctrl_serveStealReq_valid = stealServers_31_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_34_ctrl_stealReq_valid = stealServers_31_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_34_data_availableTask_ready = stealServers_31_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_34_data_qOutTask_valid = stealServers_31_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_34_data_qOutTask_bits = stealServers_31_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_35_ctrl_serveStealReq_valid = stealServers_32_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_35_ctrl_stealReq_valid = stealServers_32_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_35_data_availableTask_ready = stealServers_32_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_35_data_qOutTask_valid = stealServers_32_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_35_data_qOutTask_bits = stealServers_32_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_36_ctrl_serveStealReq_valid = stealServers_33_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_36_ctrl_stealReq_valid = stealServers_33_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_36_data_availableTask_ready = stealServers_33_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_36_data_qOutTask_valid = stealServers_33_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_36_data_qOutTask_bits = stealServers_33_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_37_ctrl_serveStealReq_valid = stealServers_34_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_37_ctrl_stealReq_valid = stealServers_34_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_37_data_availableTask_ready = stealServers_34_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_37_data_qOutTask_valid = stealServers_34_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_37_data_qOutTask_bits = stealServers_34_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_38_ctrl_serveStealReq_valid = stealServers_35_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_38_ctrl_stealReq_valid = stealServers_35_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_38_data_availableTask_ready = stealServers_35_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_38_data_qOutTask_valid = stealServers_35_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_38_data_qOutTask_bits = stealServers_35_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_39_ctrl_serveStealReq_valid = stealServers_36_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_39_ctrl_stealReq_valid = stealServers_36_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_39_data_availableTask_ready = stealServers_36_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_39_data_qOutTask_valid = stealServers_36_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_39_data_qOutTask_bits = stealServers_36_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_40_ctrl_serveStealReq_valid = stealServers_37_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_40_ctrl_stealReq_valid = stealServers_37_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_40_data_availableTask_ready = stealServers_37_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_40_data_qOutTask_valid = stealServers_37_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_40_data_qOutTask_bits = stealServers_37_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_41_ctrl_serveStealReq_valid = stealServers_38_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_41_ctrl_stealReq_valid = stealServers_38_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_41_data_availableTask_ready = stealServers_38_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_41_data_qOutTask_valid = stealServers_38_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_41_data_qOutTask_bits = stealServers_38_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_42_ctrl_serveStealReq_valid = stealServers_39_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_42_ctrl_stealReq_valid = stealServers_39_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_42_data_availableTask_ready = stealServers_39_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_42_data_qOutTask_valid = stealServers_39_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_42_data_qOutTask_bits = stealServers_39_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_43_ctrl_serveStealReq_valid = stealServers_40_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_43_ctrl_stealReq_valid = stealServers_40_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_43_data_availableTask_ready = stealServers_40_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_43_data_qOutTask_valid = stealServers_40_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_43_data_qOutTask_bits = stealServers_40_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_44_ctrl_serveStealReq_valid = stealServers_41_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_44_ctrl_stealReq_valid = stealServers_41_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_44_data_availableTask_ready = stealServers_41_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_44_data_qOutTask_valid = stealServers_41_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_44_data_qOutTask_bits = stealServers_41_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_45_ctrl_serveStealReq_valid = stealServers_42_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_45_ctrl_stealReq_valid = stealServers_42_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_45_data_availableTask_ready = stealServers_42_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_45_data_qOutTask_valid = stealServers_42_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_45_data_qOutTask_bits = stealServers_42_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_46_ctrl_serveStealReq_valid = stealServers_43_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_46_ctrl_stealReq_valid = stealServers_43_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_46_data_availableTask_ready = stealServers_43_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_46_data_qOutTask_valid = stealServers_43_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_46_data_qOutTask_bits = stealServers_43_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_47_ctrl_serveStealReq_valid = stealServers_44_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_47_ctrl_stealReq_valid = stealServers_44_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_47_data_availableTask_ready = stealServers_44_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_47_data_qOutTask_valid = stealServers_44_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_47_data_qOutTask_bits = stealServers_44_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_48_ctrl_serveStealReq_valid = stealServers_45_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_48_ctrl_stealReq_valid = stealServers_45_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_48_data_availableTask_ready = stealServers_45_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_48_data_qOutTask_valid = stealServers_45_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_48_data_qOutTask_bits = stealServers_45_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_49_ctrl_serveStealReq_valid = stealServers_46_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_49_ctrl_stealReq_valid = stealServers_46_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_49_data_availableTask_ready = stealServers_46_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_49_data_qOutTask_valid = stealServers_46_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_49_data_qOutTask_bits = stealServers_46_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_50_ctrl_serveStealReq_valid = stealServers_47_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_50_ctrl_stealReq_valid = stealServers_47_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_50_data_availableTask_ready = stealServers_47_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_50_data_qOutTask_valid = stealServers_47_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_50_data_qOutTask_bits = stealServers_47_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_51_ctrl_serveStealReq_valid = stealServers_48_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_51_ctrl_stealReq_valid = stealServers_48_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_51_data_availableTask_ready = stealServers_48_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_51_data_qOutTask_valid = stealServers_48_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_51_data_qOutTask_bits = stealServers_48_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_52_ctrl_serveStealReq_valid = stealServers_49_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_52_ctrl_stealReq_valid = stealServers_49_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_52_data_availableTask_ready = stealServers_49_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_52_data_qOutTask_valid = stealServers_49_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_52_data_qOutTask_bits = stealServers_49_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_53_ctrl_serveStealReq_valid = stealServers_50_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_53_ctrl_stealReq_valid = stealServers_50_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_53_data_availableTask_ready = stealServers_50_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_53_data_qOutTask_valid = stealServers_50_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_53_data_qOutTask_bits = stealServers_50_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_54_ctrl_serveStealReq_valid = stealServers_51_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_54_ctrl_stealReq_valid = stealServers_51_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_54_data_availableTask_ready = stealServers_51_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_54_data_qOutTask_valid = stealServers_51_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_54_data_qOutTask_bits = stealServers_51_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_55_ctrl_serveStealReq_valid = stealServers_52_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_55_ctrl_stealReq_valid = stealServers_52_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_55_data_availableTask_ready = stealServers_52_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_55_data_qOutTask_valid = stealServers_52_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_55_data_qOutTask_bits = stealServers_52_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_56_ctrl_serveStealReq_valid = stealServers_53_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_56_ctrl_stealReq_valid = stealServers_53_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_56_data_availableTask_ready = stealServers_53_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_56_data_qOutTask_valid = stealServers_53_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_56_data_qOutTask_bits = stealServers_53_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_57_ctrl_serveStealReq_valid = stealServers_54_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_57_ctrl_stealReq_valid = stealServers_54_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_57_data_availableTask_ready = stealServers_54_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_57_data_qOutTask_valid = stealServers_54_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_57_data_qOutTask_bits = stealServers_54_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_58_ctrl_serveStealReq_valid = stealServers_55_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_58_ctrl_stealReq_valid = stealServers_55_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_58_data_availableTask_ready = stealServers_55_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_58_data_qOutTask_valid = stealServers_55_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_58_data_qOutTask_bits = stealServers_55_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_59_ctrl_serveStealReq_valid = stealServers_56_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_59_ctrl_stealReq_valid = stealServers_56_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_59_data_availableTask_ready = stealServers_56_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_59_data_qOutTask_valid = stealServers_56_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_59_data_qOutTask_bits = stealServers_56_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_60_ctrl_serveStealReq_valid = stealServers_57_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_60_ctrl_stealReq_valid = stealServers_57_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_60_data_availableTask_ready = stealServers_57_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_60_data_qOutTask_valid = stealServers_57_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_60_data_qOutTask_bits = stealServers_57_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_61_ctrl_serveStealReq_valid = stealServers_58_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_61_ctrl_stealReq_valid = stealServers_58_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_61_data_availableTask_ready = stealServers_58_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_61_data_qOutTask_valid = stealServers_58_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_61_data_qOutTask_bits = stealServers_58_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_62_ctrl_serveStealReq_valid = stealServers_59_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_62_ctrl_stealReq_valid = stealServers_59_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_62_data_availableTask_ready = stealServers_59_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_62_data_qOutTask_valid = stealServers_59_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_62_data_qOutTask_bits = stealServers_59_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_63_ctrl_serveStealReq_valid = stealServers_60_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_63_ctrl_stealReq_valid = stealServers_60_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_63_data_availableTask_ready = stealServers_60_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_63_data_qOutTask_valid = stealServers_60_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_63_data_qOutTask_bits = stealServers_60_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_64_ctrl_serveStealReq_valid = stealServers_61_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_64_ctrl_stealReq_valid = stealServers_61_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_64_data_availableTask_ready = stealServers_61_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_64_data_qOutTask_valid = stealServers_61_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_64_data_qOutTask_bits = stealServers_61_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_65_ctrl_serveStealReq_valid = stealServers_62_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_65_ctrl_stealReq_valid = stealServers_62_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_65_data_availableTask_ready = stealServers_62_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_65_data_qOutTask_valid = stealServers_62_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_65_data_qOutTask_bits = stealServers_62_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_66_ctrl_serveStealReq_valid = stealServers_63_io_connNetwork_ctrl_serveStealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_66_ctrl_stealReq_valid = stealServers_63_io_connNetwork_ctrl_stealReq_valid; // @[stealNW_TQ.scala 110:44]
  assign stealNet_io_connSS_66_data_availableTask_ready = stealServers_63_io_connNetwork_data_availableTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_66_data_qOutTask_valid = stealServers_63_io_connNetwork_data_qOutTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealNet_io_connSS_66_data_qOutTask_bits = stealServers_63_io_connNetwork_data_qOutTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_0_clock = clock;
  assign stealServers_0_reset = reset;
  assign stealServers_0_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_3_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_0_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_3_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_0_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_3_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_0_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_3_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_0_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_3_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_0_io_connQ_currLength = taskQueues_0_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_0_io_connQ_push_ready = taskQueues_0_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_0_io_connQ_pop_valid = taskQueues_0_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_0_io_connQ_pop_bits = taskQueues_0_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_1_clock = clock;
  assign stealServers_1_reset = reset;
  assign stealServers_1_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_4_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_1_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_4_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_1_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_4_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_1_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_4_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_1_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_4_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_1_io_connQ_currLength = taskQueues_1_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_1_io_connQ_push_ready = taskQueues_1_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_1_io_connQ_pop_valid = taskQueues_1_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_1_io_connQ_pop_bits = taskQueues_1_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_2_clock = clock;
  assign stealServers_2_reset = reset;
  assign stealServers_2_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_5_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_2_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_5_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_2_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_5_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_2_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_5_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_2_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_5_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_2_io_connQ_currLength = taskQueues_2_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_2_io_connQ_push_ready = taskQueues_2_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_2_io_connQ_pop_valid = taskQueues_2_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_2_io_connQ_pop_bits = taskQueues_2_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_3_clock = clock;
  assign stealServers_3_reset = reset;
  assign stealServers_3_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_6_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_3_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_6_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_3_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_6_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_3_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_6_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_3_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_6_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_3_io_connQ_currLength = taskQueues_3_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_3_io_connQ_push_ready = taskQueues_3_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_3_io_connQ_pop_valid = taskQueues_3_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_3_io_connQ_pop_bits = taskQueues_3_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_4_clock = clock;
  assign stealServers_4_reset = reset;
  assign stealServers_4_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_7_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_4_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_7_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_4_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_7_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_4_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_7_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_4_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_7_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_4_io_connQ_currLength = taskQueues_4_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_4_io_connQ_push_ready = taskQueues_4_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_4_io_connQ_pop_valid = taskQueues_4_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_4_io_connQ_pop_bits = taskQueues_4_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_5_clock = clock;
  assign stealServers_5_reset = reset;
  assign stealServers_5_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_8_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_5_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_8_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_5_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_8_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_5_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_8_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_5_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_8_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_5_io_connQ_currLength = taskQueues_5_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_5_io_connQ_push_ready = taskQueues_5_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_5_io_connQ_pop_valid = taskQueues_5_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_5_io_connQ_pop_bits = taskQueues_5_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_6_clock = clock;
  assign stealServers_6_reset = reset;
  assign stealServers_6_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_9_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_6_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_9_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_6_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_9_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_6_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_9_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_6_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_9_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_6_io_connQ_currLength = taskQueues_6_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_6_io_connQ_push_ready = taskQueues_6_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_6_io_connQ_pop_valid = taskQueues_6_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_6_io_connQ_pop_bits = taskQueues_6_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_7_clock = clock;
  assign stealServers_7_reset = reset;
  assign stealServers_7_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_10_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_7_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_10_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_7_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_10_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_7_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_10_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_7_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_10_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_7_io_connQ_currLength = taskQueues_7_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_7_io_connQ_push_ready = taskQueues_7_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_7_io_connQ_pop_valid = taskQueues_7_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_7_io_connQ_pop_bits = taskQueues_7_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_8_clock = clock;
  assign stealServers_8_reset = reset;
  assign stealServers_8_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_11_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_8_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_11_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_8_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_11_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_8_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_11_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_8_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_11_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_8_io_connQ_currLength = taskQueues_8_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_8_io_connQ_push_ready = taskQueues_8_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_8_io_connQ_pop_valid = taskQueues_8_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_8_io_connQ_pop_bits = taskQueues_8_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_9_clock = clock;
  assign stealServers_9_reset = reset;
  assign stealServers_9_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_12_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_9_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_12_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_9_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_12_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_9_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_12_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_9_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_12_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_9_io_connQ_currLength = taskQueues_9_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_9_io_connQ_push_ready = taskQueues_9_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_9_io_connQ_pop_valid = taskQueues_9_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_9_io_connQ_pop_bits = taskQueues_9_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_10_clock = clock;
  assign stealServers_10_reset = reset;
  assign stealServers_10_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_13_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_10_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_13_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_10_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_13_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_10_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_13_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_10_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_13_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_10_io_connQ_currLength = taskQueues_10_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_10_io_connQ_push_ready = taskQueues_10_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_10_io_connQ_pop_valid = taskQueues_10_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_10_io_connQ_pop_bits = taskQueues_10_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_11_clock = clock;
  assign stealServers_11_reset = reset;
  assign stealServers_11_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_14_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_11_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_14_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_11_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_14_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_11_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_14_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_11_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_14_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_11_io_connQ_currLength = taskQueues_11_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_11_io_connQ_push_ready = taskQueues_11_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_11_io_connQ_pop_valid = taskQueues_11_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_11_io_connQ_pop_bits = taskQueues_11_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_12_clock = clock;
  assign stealServers_12_reset = reset;
  assign stealServers_12_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_15_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_12_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_15_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_12_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_15_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_12_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_15_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_12_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_15_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_12_io_connQ_currLength = taskQueues_12_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_12_io_connQ_push_ready = taskQueues_12_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_12_io_connQ_pop_valid = taskQueues_12_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_12_io_connQ_pop_bits = taskQueues_12_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_13_clock = clock;
  assign stealServers_13_reset = reset;
  assign stealServers_13_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_16_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_13_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_16_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_13_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_16_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_13_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_16_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_13_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_16_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_13_io_connQ_currLength = taskQueues_13_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_13_io_connQ_push_ready = taskQueues_13_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_13_io_connQ_pop_valid = taskQueues_13_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_13_io_connQ_pop_bits = taskQueues_13_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_14_clock = clock;
  assign stealServers_14_reset = reset;
  assign stealServers_14_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_17_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_14_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_17_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_14_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_17_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_14_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_17_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_14_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_17_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_14_io_connQ_currLength = taskQueues_14_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_14_io_connQ_push_ready = taskQueues_14_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_14_io_connQ_pop_valid = taskQueues_14_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_14_io_connQ_pop_bits = taskQueues_14_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_15_clock = clock;
  assign stealServers_15_reset = reset;
  assign stealServers_15_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_18_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_15_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_18_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_15_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_18_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_15_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_18_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_15_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_18_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_15_io_connQ_currLength = taskQueues_15_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_15_io_connQ_push_ready = taskQueues_15_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_15_io_connQ_pop_valid = taskQueues_15_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_15_io_connQ_pop_bits = taskQueues_15_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_16_clock = clock;
  assign stealServers_16_reset = reset;
  assign stealServers_16_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_19_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_16_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_19_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_16_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_19_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_16_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_19_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_16_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_19_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_16_io_connQ_currLength = taskQueues_16_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_16_io_connQ_push_ready = taskQueues_16_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_16_io_connQ_pop_valid = taskQueues_16_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_16_io_connQ_pop_bits = taskQueues_16_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_17_clock = clock;
  assign stealServers_17_reset = reset;
  assign stealServers_17_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_20_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_17_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_20_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_17_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_20_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_17_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_20_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_17_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_20_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_17_io_connQ_currLength = taskQueues_17_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_17_io_connQ_push_ready = taskQueues_17_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_17_io_connQ_pop_valid = taskQueues_17_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_17_io_connQ_pop_bits = taskQueues_17_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_18_clock = clock;
  assign stealServers_18_reset = reset;
  assign stealServers_18_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_21_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_18_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_21_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_18_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_21_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_18_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_21_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_18_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_21_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_18_io_connQ_currLength = taskQueues_18_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_18_io_connQ_push_ready = taskQueues_18_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_18_io_connQ_pop_valid = taskQueues_18_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_18_io_connQ_pop_bits = taskQueues_18_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_19_clock = clock;
  assign stealServers_19_reset = reset;
  assign stealServers_19_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_22_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_19_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_22_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_19_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_22_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_19_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_22_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_19_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_22_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_19_io_connQ_currLength = taskQueues_19_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_19_io_connQ_push_ready = taskQueues_19_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_19_io_connQ_pop_valid = taskQueues_19_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_19_io_connQ_pop_bits = taskQueues_19_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_20_clock = clock;
  assign stealServers_20_reset = reset;
  assign stealServers_20_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_23_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_20_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_23_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_20_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_23_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_20_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_23_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_20_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_23_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_20_io_connQ_currLength = taskQueues_20_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_20_io_connQ_push_ready = taskQueues_20_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_20_io_connQ_pop_valid = taskQueues_20_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_20_io_connQ_pop_bits = taskQueues_20_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_21_clock = clock;
  assign stealServers_21_reset = reset;
  assign stealServers_21_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_24_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_21_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_24_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_21_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_24_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_21_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_24_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_21_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_24_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_21_io_connQ_currLength = taskQueues_21_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_21_io_connQ_push_ready = taskQueues_21_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_21_io_connQ_pop_valid = taskQueues_21_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_21_io_connQ_pop_bits = taskQueues_21_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_22_clock = clock;
  assign stealServers_22_reset = reset;
  assign stealServers_22_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_25_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_22_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_25_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_22_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_25_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_22_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_25_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_22_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_25_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_22_io_connQ_currLength = taskQueues_22_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_22_io_connQ_push_ready = taskQueues_22_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_22_io_connQ_pop_valid = taskQueues_22_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_22_io_connQ_pop_bits = taskQueues_22_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_23_clock = clock;
  assign stealServers_23_reset = reset;
  assign stealServers_23_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_26_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_23_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_26_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_23_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_26_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_23_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_26_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_23_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_26_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_23_io_connQ_currLength = taskQueues_23_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_23_io_connQ_push_ready = taskQueues_23_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_23_io_connQ_pop_valid = taskQueues_23_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_23_io_connQ_pop_bits = taskQueues_23_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_24_clock = clock;
  assign stealServers_24_reset = reset;
  assign stealServers_24_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_27_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_24_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_27_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_24_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_27_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_24_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_27_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_24_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_27_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_24_io_connQ_currLength = taskQueues_24_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_24_io_connQ_push_ready = taskQueues_24_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_24_io_connQ_pop_valid = taskQueues_24_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_24_io_connQ_pop_bits = taskQueues_24_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_25_clock = clock;
  assign stealServers_25_reset = reset;
  assign stealServers_25_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_28_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_25_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_28_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_25_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_28_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_25_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_28_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_25_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_28_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_25_io_connQ_currLength = taskQueues_25_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_25_io_connQ_push_ready = taskQueues_25_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_25_io_connQ_pop_valid = taskQueues_25_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_25_io_connQ_pop_bits = taskQueues_25_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_26_clock = clock;
  assign stealServers_26_reset = reset;
  assign stealServers_26_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_29_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_26_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_29_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_26_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_29_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_26_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_29_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_26_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_29_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_26_io_connQ_currLength = taskQueues_26_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_26_io_connQ_push_ready = taskQueues_26_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_26_io_connQ_pop_valid = taskQueues_26_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_26_io_connQ_pop_bits = taskQueues_26_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_27_clock = clock;
  assign stealServers_27_reset = reset;
  assign stealServers_27_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_30_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_27_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_30_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_27_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_30_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_27_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_30_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_27_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_30_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_27_io_connQ_currLength = taskQueues_27_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_27_io_connQ_push_ready = taskQueues_27_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_27_io_connQ_pop_valid = taskQueues_27_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_27_io_connQ_pop_bits = taskQueues_27_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_28_clock = clock;
  assign stealServers_28_reset = reset;
  assign stealServers_28_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_31_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_28_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_31_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_28_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_31_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_28_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_31_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_28_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_31_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_28_io_connQ_currLength = taskQueues_28_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_28_io_connQ_push_ready = taskQueues_28_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_28_io_connQ_pop_valid = taskQueues_28_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_28_io_connQ_pop_bits = taskQueues_28_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_29_clock = clock;
  assign stealServers_29_reset = reset;
  assign stealServers_29_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_32_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_29_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_32_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_29_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_32_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_29_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_32_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_29_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_32_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_29_io_connQ_currLength = taskQueues_29_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_29_io_connQ_push_ready = taskQueues_29_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_29_io_connQ_pop_valid = taskQueues_29_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_29_io_connQ_pop_bits = taskQueues_29_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_30_clock = clock;
  assign stealServers_30_reset = reset;
  assign stealServers_30_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_33_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_30_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_33_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_30_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_33_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_30_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_33_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_30_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_33_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_30_io_connQ_currLength = taskQueues_30_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_30_io_connQ_push_ready = taskQueues_30_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_30_io_connQ_pop_valid = taskQueues_30_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_30_io_connQ_pop_bits = taskQueues_30_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_31_clock = clock;
  assign stealServers_31_reset = reset;
  assign stealServers_31_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_34_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_31_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_34_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_31_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_34_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_31_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_34_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_31_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_34_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_31_io_connQ_currLength = taskQueues_31_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_31_io_connQ_push_ready = taskQueues_31_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_31_io_connQ_pop_valid = taskQueues_31_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_31_io_connQ_pop_bits = taskQueues_31_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_32_clock = clock;
  assign stealServers_32_reset = reset;
  assign stealServers_32_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_35_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_32_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_35_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_32_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_35_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_32_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_35_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_32_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_35_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_32_io_connQ_currLength = taskQueues_32_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_32_io_connQ_push_ready = taskQueues_32_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_32_io_connQ_pop_valid = taskQueues_32_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_32_io_connQ_pop_bits = taskQueues_32_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_33_clock = clock;
  assign stealServers_33_reset = reset;
  assign stealServers_33_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_36_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_33_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_36_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_33_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_36_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_33_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_36_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_33_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_36_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_33_io_connQ_currLength = taskQueues_33_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_33_io_connQ_push_ready = taskQueues_33_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_33_io_connQ_pop_valid = taskQueues_33_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_33_io_connQ_pop_bits = taskQueues_33_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_34_clock = clock;
  assign stealServers_34_reset = reset;
  assign stealServers_34_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_37_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_34_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_37_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_34_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_37_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_34_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_37_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_34_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_37_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_34_io_connQ_currLength = taskQueues_34_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_34_io_connQ_push_ready = taskQueues_34_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_34_io_connQ_pop_valid = taskQueues_34_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_34_io_connQ_pop_bits = taskQueues_34_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_35_clock = clock;
  assign stealServers_35_reset = reset;
  assign stealServers_35_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_38_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_35_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_38_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_35_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_38_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_35_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_38_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_35_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_38_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_35_io_connQ_currLength = taskQueues_35_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_35_io_connQ_push_ready = taskQueues_35_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_35_io_connQ_pop_valid = taskQueues_35_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_35_io_connQ_pop_bits = taskQueues_35_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_36_clock = clock;
  assign stealServers_36_reset = reset;
  assign stealServers_36_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_39_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_36_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_39_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_36_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_39_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_36_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_39_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_36_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_39_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_36_io_connQ_currLength = taskQueues_36_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_36_io_connQ_push_ready = taskQueues_36_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_36_io_connQ_pop_valid = taskQueues_36_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_36_io_connQ_pop_bits = taskQueues_36_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_37_clock = clock;
  assign stealServers_37_reset = reset;
  assign stealServers_37_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_40_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_37_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_40_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_37_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_40_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_37_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_40_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_37_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_40_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_37_io_connQ_currLength = taskQueues_37_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_37_io_connQ_push_ready = taskQueues_37_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_37_io_connQ_pop_valid = taskQueues_37_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_37_io_connQ_pop_bits = taskQueues_37_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_38_clock = clock;
  assign stealServers_38_reset = reset;
  assign stealServers_38_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_41_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_38_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_41_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_38_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_41_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_38_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_41_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_38_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_41_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_38_io_connQ_currLength = taskQueues_38_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_38_io_connQ_push_ready = taskQueues_38_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_38_io_connQ_pop_valid = taskQueues_38_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_38_io_connQ_pop_bits = taskQueues_38_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_39_clock = clock;
  assign stealServers_39_reset = reset;
  assign stealServers_39_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_42_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_39_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_42_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_39_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_42_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_39_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_42_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_39_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_42_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_39_io_connQ_currLength = taskQueues_39_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_39_io_connQ_push_ready = taskQueues_39_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_39_io_connQ_pop_valid = taskQueues_39_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_39_io_connQ_pop_bits = taskQueues_39_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_40_clock = clock;
  assign stealServers_40_reset = reset;
  assign stealServers_40_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_43_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_40_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_43_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_40_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_43_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_40_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_43_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_40_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_43_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_40_io_connQ_currLength = taskQueues_40_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_40_io_connQ_push_ready = taskQueues_40_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_40_io_connQ_pop_valid = taskQueues_40_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_40_io_connQ_pop_bits = taskQueues_40_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_41_clock = clock;
  assign stealServers_41_reset = reset;
  assign stealServers_41_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_44_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_41_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_44_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_41_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_44_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_41_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_44_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_41_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_44_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_41_io_connQ_currLength = taskQueues_41_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_41_io_connQ_push_ready = taskQueues_41_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_41_io_connQ_pop_valid = taskQueues_41_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_41_io_connQ_pop_bits = taskQueues_41_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_42_clock = clock;
  assign stealServers_42_reset = reset;
  assign stealServers_42_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_45_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_42_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_45_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_42_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_45_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_42_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_45_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_42_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_45_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_42_io_connQ_currLength = taskQueues_42_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_42_io_connQ_push_ready = taskQueues_42_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_42_io_connQ_pop_valid = taskQueues_42_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_42_io_connQ_pop_bits = taskQueues_42_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_43_clock = clock;
  assign stealServers_43_reset = reset;
  assign stealServers_43_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_46_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_43_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_46_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_43_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_46_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_43_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_46_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_43_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_46_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_43_io_connQ_currLength = taskQueues_43_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_43_io_connQ_push_ready = taskQueues_43_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_43_io_connQ_pop_valid = taskQueues_43_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_43_io_connQ_pop_bits = taskQueues_43_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_44_clock = clock;
  assign stealServers_44_reset = reset;
  assign stealServers_44_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_47_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_44_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_47_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_44_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_47_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_44_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_47_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_44_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_47_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_44_io_connQ_currLength = taskQueues_44_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_44_io_connQ_push_ready = taskQueues_44_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_44_io_connQ_pop_valid = taskQueues_44_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_44_io_connQ_pop_bits = taskQueues_44_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_45_clock = clock;
  assign stealServers_45_reset = reset;
  assign stealServers_45_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_48_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_45_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_48_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_45_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_48_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_45_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_48_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_45_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_48_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_45_io_connQ_currLength = taskQueues_45_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_45_io_connQ_push_ready = taskQueues_45_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_45_io_connQ_pop_valid = taskQueues_45_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_45_io_connQ_pop_bits = taskQueues_45_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_46_clock = clock;
  assign stealServers_46_reset = reset;
  assign stealServers_46_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_49_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_46_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_49_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_46_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_49_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_46_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_49_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_46_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_49_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_46_io_connQ_currLength = taskQueues_46_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_46_io_connQ_push_ready = taskQueues_46_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_46_io_connQ_pop_valid = taskQueues_46_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_46_io_connQ_pop_bits = taskQueues_46_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_47_clock = clock;
  assign stealServers_47_reset = reset;
  assign stealServers_47_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_50_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_47_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_50_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_47_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_50_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_47_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_50_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_47_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_50_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_47_io_connQ_currLength = taskQueues_47_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_47_io_connQ_push_ready = taskQueues_47_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_47_io_connQ_pop_valid = taskQueues_47_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_47_io_connQ_pop_bits = taskQueues_47_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_48_clock = clock;
  assign stealServers_48_reset = reset;
  assign stealServers_48_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_51_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_48_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_51_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_48_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_51_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_48_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_51_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_48_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_51_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_48_io_connQ_currLength = taskQueues_48_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_48_io_connQ_push_ready = taskQueues_48_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_48_io_connQ_pop_valid = taskQueues_48_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_48_io_connQ_pop_bits = taskQueues_48_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_49_clock = clock;
  assign stealServers_49_reset = reset;
  assign stealServers_49_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_52_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_49_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_52_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_49_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_52_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_49_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_52_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_49_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_52_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_49_io_connQ_currLength = taskQueues_49_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_49_io_connQ_push_ready = taskQueues_49_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_49_io_connQ_pop_valid = taskQueues_49_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_49_io_connQ_pop_bits = taskQueues_49_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_50_clock = clock;
  assign stealServers_50_reset = reset;
  assign stealServers_50_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_53_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_50_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_53_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_50_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_53_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_50_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_53_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_50_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_53_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_50_io_connQ_currLength = taskQueues_50_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_50_io_connQ_push_ready = taskQueues_50_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_50_io_connQ_pop_valid = taskQueues_50_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_50_io_connQ_pop_bits = taskQueues_50_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_51_clock = clock;
  assign stealServers_51_reset = reset;
  assign stealServers_51_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_54_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_51_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_54_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_51_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_54_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_51_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_54_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_51_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_54_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_51_io_connQ_currLength = taskQueues_51_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_51_io_connQ_push_ready = taskQueues_51_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_51_io_connQ_pop_valid = taskQueues_51_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_51_io_connQ_pop_bits = taskQueues_51_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_52_clock = clock;
  assign stealServers_52_reset = reset;
  assign stealServers_52_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_55_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_52_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_55_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_52_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_55_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_52_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_55_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_52_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_55_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_52_io_connQ_currLength = taskQueues_52_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_52_io_connQ_push_ready = taskQueues_52_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_52_io_connQ_pop_valid = taskQueues_52_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_52_io_connQ_pop_bits = taskQueues_52_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_53_clock = clock;
  assign stealServers_53_reset = reset;
  assign stealServers_53_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_56_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_53_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_56_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_53_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_56_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_53_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_56_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_53_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_56_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_53_io_connQ_currLength = taskQueues_53_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_53_io_connQ_push_ready = taskQueues_53_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_53_io_connQ_pop_valid = taskQueues_53_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_53_io_connQ_pop_bits = taskQueues_53_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_54_clock = clock;
  assign stealServers_54_reset = reset;
  assign stealServers_54_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_57_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_54_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_57_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_54_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_57_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_54_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_57_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_54_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_57_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_54_io_connQ_currLength = taskQueues_54_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_54_io_connQ_push_ready = taskQueues_54_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_54_io_connQ_pop_valid = taskQueues_54_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_54_io_connQ_pop_bits = taskQueues_54_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_55_clock = clock;
  assign stealServers_55_reset = reset;
  assign stealServers_55_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_58_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_55_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_58_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_55_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_58_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_55_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_58_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_55_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_58_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_55_io_connQ_currLength = taskQueues_55_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_55_io_connQ_push_ready = taskQueues_55_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_55_io_connQ_pop_valid = taskQueues_55_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_55_io_connQ_pop_bits = taskQueues_55_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_56_clock = clock;
  assign stealServers_56_reset = reset;
  assign stealServers_56_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_59_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_56_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_59_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_56_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_59_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_56_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_59_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_56_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_59_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_56_io_connQ_currLength = taskQueues_56_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_56_io_connQ_push_ready = taskQueues_56_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_56_io_connQ_pop_valid = taskQueues_56_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_56_io_connQ_pop_bits = taskQueues_56_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_57_clock = clock;
  assign stealServers_57_reset = reset;
  assign stealServers_57_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_60_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_57_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_60_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_57_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_60_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_57_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_60_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_57_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_60_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_57_io_connQ_currLength = taskQueues_57_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_57_io_connQ_push_ready = taskQueues_57_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_57_io_connQ_pop_valid = taskQueues_57_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_57_io_connQ_pop_bits = taskQueues_57_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_58_clock = clock;
  assign stealServers_58_reset = reset;
  assign stealServers_58_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_61_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_58_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_61_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_58_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_61_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_58_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_61_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_58_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_61_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_58_io_connQ_currLength = taskQueues_58_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_58_io_connQ_push_ready = taskQueues_58_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_58_io_connQ_pop_valid = taskQueues_58_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_58_io_connQ_pop_bits = taskQueues_58_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_59_clock = clock;
  assign stealServers_59_reset = reset;
  assign stealServers_59_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_62_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_59_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_62_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_59_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_62_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_59_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_62_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_59_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_62_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_59_io_connQ_currLength = taskQueues_59_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_59_io_connQ_push_ready = taskQueues_59_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_59_io_connQ_pop_valid = taskQueues_59_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_59_io_connQ_pop_bits = taskQueues_59_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_60_clock = clock;
  assign stealServers_60_reset = reset;
  assign stealServers_60_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_63_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_60_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_63_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_60_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_63_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_60_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_63_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_60_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_63_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_60_io_connQ_currLength = taskQueues_60_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_60_io_connQ_push_ready = taskQueues_60_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_60_io_connQ_pop_valid = taskQueues_60_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_60_io_connQ_pop_bits = taskQueues_60_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_61_clock = clock;
  assign stealServers_61_reset = reset;
  assign stealServers_61_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_64_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_61_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_64_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_61_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_64_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_61_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_64_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_61_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_64_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_61_io_connQ_currLength = taskQueues_61_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_61_io_connQ_push_ready = taskQueues_61_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_61_io_connQ_pop_valid = taskQueues_61_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_61_io_connQ_pop_bits = taskQueues_61_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_62_clock = clock;
  assign stealServers_62_reset = reset;
  assign stealServers_62_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_65_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_62_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_65_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_62_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_65_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_62_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_65_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_62_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_65_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_62_io_connQ_currLength = taskQueues_62_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_62_io_connQ_push_ready = taskQueues_62_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_62_io_connQ_pop_valid = taskQueues_62_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_62_io_connQ_pop_bits = taskQueues_62_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign stealServers_63_clock = clock;
  assign stealServers_63_reset = reset;
  assign stealServers_63_io_connNetwork_ctrl_serveStealReq_ready = stealNet_io_connSS_66_ctrl_serveStealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_63_io_connNetwork_ctrl_stealReq_ready = stealNet_io_connSS_66_ctrl_stealReq_ready; // @[stealNW_TQ.scala 110:44]
  assign stealServers_63_io_connNetwork_data_availableTask_valid = stealNet_io_connSS_66_data_availableTask_valid; // @[stealNW_TQ.scala 93:44]
  assign stealServers_63_io_connNetwork_data_availableTask_bits = stealNet_io_connSS_66_data_availableTask_bits; // @[stealNW_TQ.scala 93:44]
  assign stealServers_63_io_connNetwork_data_qOutTask_ready = stealNet_io_connSS_66_data_qOutTask_ready; // @[stealNW_TQ.scala 93:44]
  assign stealServers_63_io_connQ_currLength = taskQueues_63_io_connVec_1_currLength[5:0]; // @[stealNW_TQ.scala 69:37]
  assign stealServers_63_io_connQ_push_ready = taskQueues_63_io_connVec_1_push_ready; // @[stealNW_TQ.scala 69:37]
  assign stealServers_63_io_connQ_pop_valid = taskQueues_63_io_connVec_1_pop_valid; // @[stealNW_TQ.scala 69:37]
  assign stealServers_63_io_connQ_pop_bits = taskQueues_63_io_connVec_1_pop_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_0_clock = clock;
  assign taskQueues_0_reset = reset;
  assign taskQueues_0_io_connVec_0_push_valid = io_connPE_0_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_0_io_connVec_0_push_bits = io_connPE_0_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_0_io_connVec_0_pop_ready = io_connPE_0_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_0_io_connVec_1_push_valid = stealServers_0_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_0_io_connVec_1_push_bits = stealServers_0_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_0_io_connVec_1_pop_ready = stealServers_0_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_1_clock = clock;
  assign taskQueues_1_reset = reset;
  assign taskQueues_1_io_connVec_0_push_valid = io_connPE_1_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_1_io_connVec_0_push_bits = io_connPE_1_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_1_io_connVec_0_pop_ready = io_connPE_1_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_1_io_connVec_1_push_valid = stealServers_1_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_1_io_connVec_1_push_bits = stealServers_1_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_1_io_connVec_1_pop_ready = stealServers_1_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_2_clock = clock;
  assign taskQueues_2_reset = reset;
  assign taskQueues_2_io_connVec_0_push_valid = io_connPE_2_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_2_io_connVec_0_push_bits = io_connPE_2_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_2_io_connVec_0_pop_ready = io_connPE_2_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_2_io_connVec_1_push_valid = stealServers_2_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_2_io_connVec_1_push_bits = stealServers_2_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_2_io_connVec_1_pop_ready = stealServers_2_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_3_clock = clock;
  assign taskQueues_3_reset = reset;
  assign taskQueues_3_io_connVec_0_push_valid = io_connPE_3_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_3_io_connVec_0_push_bits = io_connPE_3_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_3_io_connVec_0_pop_ready = io_connPE_3_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_3_io_connVec_1_push_valid = stealServers_3_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_3_io_connVec_1_push_bits = stealServers_3_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_3_io_connVec_1_pop_ready = stealServers_3_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_4_clock = clock;
  assign taskQueues_4_reset = reset;
  assign taskQueues_4_io_connVec_0_push_valid = io_connPE_4_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_4_io_connVec_0_push_bits = io_connPE_4_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_4_io_connVec_0_pop_ready = io_connPE_4_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_4_io_connVec_1_push_valid = stealServers_4_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_4_io_connVec_1_push_bits = stealServers_4_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_4_io_connVec_1_pop_ready = stealServers_4_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_5_clock = clock;
  assign taskQueues_5_reset = reset;
  assign taskQueues_5_io_connVec_0_push_valid = io_connPE_5_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_5_io_connVec_0_push_bits = io_connPE_5_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_5_io_connVec_0_pop_ready = io_connPE_5_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_5_io_connVec_1_push_valid = stealServers_5_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_5_io_connVec_1_push_bits = stealServers_5_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_5_io_connVec_1_pop_ready = stealServers_5_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_6_clock = clock;
  assign taskQueues_6_reset = reset;
  assign taskQueues_6_io_connVec_0_push_valid = io_connPE_6_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_6_io_connVec_0_push_bits = io_connPE_6_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_6_io_connVec_0_pop_ready = io_connPE_6_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_6_io_connVec_1_push_valid = stealServers_6_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_6_io_connVec_1_push_bits = stealServers_6_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_6_io_connVec_1_pop_ready = stealServers_6_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_7_clock = clock;
  assign taskQueues_7_reset = reset;
  assign taskQueues_7_io_connVec_0_push_valid = io_connPE_7_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_7_io_connVec_0_push_bits = io_connPE_7_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_7_io_connVec_0_pop_ready = io_connPE_7_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_7_io_connVec_1_push_valid = stealServers_7_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_7_io_connVec_1_push_bits = stealServers_7_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_7_io_connVec_1_pop_ready = stealServers_7_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_8_clock = clock;
  assign taskQueues_8_reset = reset;
  assign taskQueues_8_io_connVec_0_push_valid = io_connPE_8_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_8_io_connVec_0_push_bits = io_connPE_8_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_8_io_connVec_0_pop_ready = io_connPE_8_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_8_io_connVec_1_push_valid = stealServers_8_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_8_io_connVec_1_push_bits = stealServers_8_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_8_io_connVec_1_pop_ready = stealServers_8_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_9_clock = clock;
  assign taskQueues_9_reset = reset;
  assign taskQueues_9_io_connVec_0_push_valid = io_connPE_9_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_9_io_connVec_0_push_bits = io_connPE_9_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_9_io_connVec_0_pop_ready = io_connPE_9_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_9_io_connVec_1_push_valid = stealServers_9_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_9_io_connVec_1_push_bits = stealServers_9_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_9_io_connVec_1_pop_ready = stealServers_9_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_10_clock = clock;
  assign taskQueues_10_reset = reset;
  assign taskQueues_10_io_connVec_0_push_valid = io_connPE_10_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_10_io_connVec_0_push_bits = io_connPE_10_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_10_io_connVec_0_pop_ready = io_connPE_10_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_10_io_connVec_1_push_valid = stealServers_10_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_10_io_connVec_1_push_bits = stealServers_10_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_10_io_connVec_1_pop_ready = stealServers_10_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_11_clock = clock;
  assign taskQueues_11_reset = reset;
  assign taskQueues_11_io_connVec_0_push_valid = io_connPE_11_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_11_io_connVec_0_push_bits = io_connPE_11_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_11_io_connVec_0_pop_ready = io_connPE_11_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_11_io_connVec_1_push_valid = stealServers_11_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_11_io_connVec_1_push_bits = stealServers_11_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_11_io_connVec_1_pop_ready = stealServers_11_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_12_clock = clock;
  assign taskQueues_12_reset = reset;
  assign taskQueues_12_io_connVec_0_push_valid = io_connPE_12_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_12_io_connVec_0_push_bits = io_connPE_12_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_12_io_connVec_0_pop_ready = io_connPE_12_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_12_io_connVec_1_push_valid = stealServers_12_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_12_io_connVec_1_push_bits = stealServers_12_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_12_io_connVec_1_pop_ready = stealServers_12_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_13_clock = clock;
  assign taskQueues_13_reset = reset;
  assign taskQueues_13_io_connVec_0_push_valid = io_connPE_13_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_13_io_connVec_0_push_bits = io_connPE_13_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_13_io_connVec_0_pop_ready = io_connPE_13_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_13_io_connVec_1_push_valid = stealServers_13_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_13_io_connVec_1_push_bits = stealServers_13_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_13_io_connVec_1_pop_ready = stealServers_13_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_14_clock = clock;
  assign taskQueues_14_reset = reset;
  assign taskQueues_14_io_connVec_0_push_valid = io_connPE_14_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_14_io_connVec_0_push_bits = io_connPE_14_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_14_io_connVec_0_pop_ready = io_connPE_14_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_14_io_connVec_1_push_valid = stealServers_14_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_14_io_connVec_1_push_bits = stealServers_14_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_14_io_connVec_1_pop_ready = stealServers_14_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_15_clock = clock;
  assign taskQueues_15_reset = reset;
  assign taskQueues_15_io_connVec_0_push_valid = io_connPE_15_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_15_io_connVec_0_push_bits = io_connPE_15_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_15_io_connVec_0_pop_ready = io_connPE_15_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_15_io_connVec_1_push_valid = stealServers_15_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_15_io_connVec_1_push_bits = stealServers_15_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_15_io_connVec_1_pop_ready = stealServers_15_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_16_clock = clock;
  assign taskQueues_16_reset = reset;
  assign taskQueues_16_io_connVec_0_push_valid = io_connPE_16_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_16_io_connVec_0_push_bits = io_connPE_16_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_16_io_connVec_0_pop_ready = io_connPE_16_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_16_io_connVec_1_push_valid = stealServers_16_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_16_io_connVec_1_push_bits = stealServers_16_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_16_io_connVec_1_pop_ready = stealServers_16_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_17_clock = clock;
  assign taskQueues_17_reset = reset;
  assign taskQueues_17_io_connVec_0_push_valid = io_connPE_17_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_17_io_connVec_0_push_bits = io_connPE_17_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_17_io_connVec_0_pop_ready = io_connPE_17_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_17_io_connVec_1_push_valid = stealServers_17_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_17_io_connVec_1_push_bits = stealServers_17_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_17_io_connVec_1_pop_ready = stealServers_17_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_18_clock = clock;
  assign taskQueues_18_reset = reset;
  assign taskQueues_18_io_connVec_0_push_valid = io_connPE_18_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_18_io_connVec_0_push_bits = io_connPE_18_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_18_io_connVec_0_pop_ready = io_connPE_18_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_18_io_connVec_1_push_valid = stealServers_18_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_18_io_connVec_1_push_bits = stealServers_18_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_18_io_connVec_1_pop_ready = stealServers_18_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_19_clock = clock;
  assign taskQueues_19_reset = reset;
  assign taskQueues_19_io_connVec_0_push_valid = io_connPE_19_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_19_io_connVec_0_push_bits = io_connPE_19_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_19_io_connVec_0_pop_ready = io_connPE_19_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_19_io_connVec_1_push_valid = stealServers_19_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_19_io_connVec_1_push_bits = stealServers_19_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_19_io_connVec_1_pop_ready = stealServers_19_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_20_clock = clock;
  assign taskQueues_20_reset = reset;
  assign taskQueues_20_io_connVec_0_push_valid = io_connPE_20_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_20_io_connVec_0_push_bits = io_connPE_20_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_20_io_connVec_0_pop_ready = io_connPE_20_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_20_io_connVec_1_push_valid = stealServers_20_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_20_io_connVec_1_push_bits = stealServers_20_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_20_io_connVec_1_pop_ready = stealServers_20_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_21_clock = clock;
  assign taskQueues_21_reset = reset;
  assign taskQueues_21_io_connVec_0_push_valid = io_connPE_21_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_21_io_connVec_0_push_bits = io_connPE_21_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_21_io_connVec_0_pop_ready = io_connPE_21_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_21_io_connVec_1_push_valid = stealServers_21_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_21_io_connVec_1_push_bits = stealServers_21_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_21_io_connVec_1_pop_ready = stealServers_21_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_22_clock = clock;
  assign taskQueues_22_reset = reset;
  assign taskQueues_22_io_connVec_0_push_valid = io_connPE_22_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_22_io_connVec_0_push_bits = io_connPE_22_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_22_io_connVec_0_pop_ready = io_connPE_22_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_22_io_connVec_1_push_valid = stealServers_22_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_22_io_connVec_1_push_bits = stealServers_22_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_22_io_connVec_1_pop_ready = stealServers_22_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_23_clock = clock;
  assign taskQueues_23_reset = reset;
  assign taskQueues_23_io_connVec_0_push_valid = io_connPE_23_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_23_io_connVec_0_push_bits = io_connPE_23_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_23_io_connVec_0_pop_ready = io_connPE_23_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_23_io_connVec_1_push_valid = stealServers_23_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_23_io_connVec_1_push_bits = stealServers_23_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_23_io_connVec_1_pop_ready = stealServers_23_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_24_clock = clock;
  assign taskQueues_24_reset = reset;
  assign taskQueues_24_io_connVec_0_push_valid = io_connPE_24_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_24_io_connVec_0_push_bits = io_connPE_24_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_24_io_connVec_0_pop_ready = io_connPE_24_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_24_io_connVec_1_push_valid = stealServers_24_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_24_io_connVec_1_push_bits = stealServers_24_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_24_io_connVec_1_pop_ready = stealServers_24_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_25_clock = clock;
  assign taskQueues_25_reset = reset;
  assign taskQueues_25_io_connVec_0_push_valid = io_connPE_25_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_25_io_connVec_0_push_bits = io_connPE_25_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_25_io_connVec_0_pop_ready = io_connPE_25_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_25_io_connVec_1_push_valid = stealServers_25_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_25_io_connVec_1_push_bits = stealServers_25_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_25_io_connVec_1_pop_ready = stealServers_25_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_26_clock = clock;
  assign taskQueues_26_reset = reset;
  assign taskQueues_26_io_connVec_0_push_valid = io_connPE_26_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_26_io_connVec_0_push_bits = io_connPE_26_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_26_io_connVec_0_pop_ready = io_connPE_26_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_26_io_connVec_1_push_valid = stealServers_26_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_26_io_connVec_1_push_bits = stealServers_26_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_26_io_connVec_1_pop_ready = stealServers_26_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_27_clock = clock;
  assign taskQueues_27_reset = reset;
  assign taskQueues_27_io_connVec_0_push_valid = io_connPE_27_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_27_io_connVec_0_push_bits = io_connPE_27_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_27_io_connVec_0_pop_ready = io_connPE_27_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_27_io_connVec_1_push_valid = stealServers_27_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_27_io_connVec_1_push_bits = stealServers_27_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_27_io_connVec_1_pop_ready = stealServers_27_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_28_clock = clock;
  assign taskQueues_28_reset = reset;
  assign taskQueues_28_io_connVec_0_push_valid = io_connPE_28_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_28_io_connVec_0_push_bits = io_connPE_28_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_28_io_connVec_0_pop_ready = io_connPE_28_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_28_io_connVec_1_push_valid = stealServers_28_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_28_io_connVec_1_push_bits = stealServers_28_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_28_io_connVec_1_pop_ready = stealServers_28_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_29_clock = clock;
  assign taskQueues_29_reset = reset;
  assign taskQueues_29_io_connVec_0_push_valid = io_connPE_29_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_29_io_connVec_0_push_bits = io_connPE_29_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_29_io_connVec_0_pop_ready = io_connPE_29_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_29_io_connVec_1_push_valid = stealServers_29_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_29_io_connVec_1_push_bits = stealServers_29_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_29_io_connVec_1_pop_ready = stealServers_29_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_30_clock = clock;
  assign taskQueues_30_reset = reset;
  assign taskQueues_30_io_connVec_0_push_valid = io_connPE_30_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_30_io_connVec_0_push_bits = io_connPE_30_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_30_io_connVec_0_pop_ready = io_connPE_30_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_30_io_connVec_1_push_valid = stealServers_30_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_30_io_connVec_1_push_bits = stealServers_30_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_30_io_connVec_1_pop_ready = stealServers_30_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_31_clock = clock;
  assign taskQueues_31_reset = reset;
  assign taskQueues_31_io_connVec_0_push_valid = io_connPE_31_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_31_io_connVec_0_push_bits = io_connPE_31_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_31_io_connVec_0_pop_ready = io_connPE_31_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_31_io_connVec_1_push_valid = stealServers_31_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_31_io_connVec_1_push_bits = stealServers_31_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_31_io_connVec_1_pop_ready = stealServers_31_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_32_clock = clock;
  assign taskQueues_32_reset = reset;
  assign taskQueues_32_io_connVec_0_push_valid = io_connPE_32_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_32_io_connVec_0_push_bits = io_connPE_32_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_32_io_connVec_0_pop_ready = io_connPE_32_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_32_io_connVec_1_push_valid = stealServers_32_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_32_io_connVec_1_push_bits = stealServers_32_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_32_io_connVec_1_pop_ready = stealServers_32_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_33_clock = clock;
  assign taskQueues_33_reset = reset;
  assign taskQueues_33_io_connVec_0_push_valid = io_connPE_33_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_33_io_connVec_0_push_bits = io_connPE_33_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_33_io_connVec_0_pop_ready = io_connPE_33_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_33_io_connVec_1_push_valid = stealServers_33_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_33_io_connVec_1_push_bits = stealServers_33_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_33_io_connVec_1_pop_ready = stealServers_33_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_34_clock = clock;
  assign taskQueues_34_reset = reset;
  assign taskQueues_34_io_connVec_0_push_valid = io_connPE_34_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_34_io_connVec_0_push_bits = io_connPE_34_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_34_io_connVec_0_pop_ready = io_connPE_34_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_34_io_connVec_1_push_valid = stealServers_34_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_34_io_connVec_1_push_bits = stealServers_34_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_34_io_connVec_1_pop_ready = stealServers_34_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_35_clock = clock;
  assign taskQueues_35_reset = reset;
  assign taskQueues_35_io_connVec_0_push_valid = io_connPE_35_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_35_io_connVec_0_push_bits = io_connPE_35_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_35_io_connVec_0_pop_ready = io_connPE_35_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_35_io_connVec_1_push_valid = stealServers_35_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_35_io_connVec_1_push_bits = stealServers_35_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_35_io_connVec_1_pop_ready = stealServers_35_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_36_clock = clock;
  assign taskQueues_36_reset = reset;
  assign taskQueues_36_io_connVec_0_push_valid = io_connPE_36_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_36_io_connVec_0_push_bits = io_connPE_36_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_36_io_connVec_0_pop_ready = io_connPE_36_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_36_io_connVec_1_push_valid = stealServers_36_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_36_io_connVec_1_push_bits = stealServers_36_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_36_io_connVec_1_pop_ready = stealServers_36_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_37_clock = clock;
  assign taskQueues_37_reset = reset;
  assign taskQueues_37_io_connVec_0_push_valid = io_connPE_37_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_37_io_connVec_0_push_bits = io_connPE_37_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_37_io_connVec_0_pop_ready = io_connPE_37_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_37_io_connVec_1_push_valid = stealServers_37_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_37_io_connVec_1_push_bits = stealServers_37_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_37_io_connVec_1_pop_ready = stealServers_37_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_38_clock = clock;
  assign taskQueues_38_reset = reset;
  assign taskQueues_38_io_connVec_0_push_valid = io_connPE_38_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_38_io_connVec_0_push_bits = io_connPE_38_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_38_io_connVec_0_pop_ready = io_connPE_38_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_38_io_connVec_1_push_valid = stealServers_38_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_38_io_connVec_1_push_bits = stealServers_38_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_38_io_connVec_1_pop_ready = stealServers_38_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_39_clock = clock;
  assign taskQueues_39_reset = reset;
  assign taskQueues_39_io_connVec_0_push_valid = io_connPE_39_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_39_io_connVec_0_push_bits = io_connPE_39_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_39_io_connVec_0_pop_ready = io_connPE_39_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_39_io_connVec_1_push_valid = stealServers_39_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_39_io_connVec_1_push_bits = stealServers_39_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_39_io_connVec_1_pop_ready = stealServers_39_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_40_clock = clock;
  assign taskQueues_40_reset = reset;
  assign taskQueues_40_io_connVec_0_push_valid = io_connPE_40_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_40_io_connVec_0_push_bits = io_connPE_40_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_40_io_connVec_0_pop_ready = io_connPE_40_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_40_io_connVec_1_push_valid = stealServers_40_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_40_io_connVec_1_push_bits = stealServers_40_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_40_io_connVec_1_pop_ready = stealServers_40_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_41_clock = clock;
  assign taskQueues_41_reset = reset;
  assign taskQueues_41_io_connVec_0_push_valid = io_connPE_41_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_41_io_connVec_0_push_bits = io_connPE_41_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_41_io_connVec_0_pop_ready = io_connPE_41_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_41_io_connVec_1_push_valid = stealServers_41_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_41_io_connVec_1_push_bits = stealServers_41_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_41_io_connVec_1_pop_ready = stealServers_41_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_42_clock = clock;
  assign taskQueues_42_reset = reset;
  assign taskQueues_42_io_connVec_0_push_valid = io_connPE_42_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_42_io_connVec_0_push_bits = io_connPE_42_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_42_io_connVec_0_pop_ready = io_connPE_42_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_42_io_connVec_1_push_valid = stealServers_42_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_42_io_connVec_1_push_bits = stealServers_42_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_42_io_connVec_1_pop_ready = stealServers_42_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_43_clock = clock;
  assign taskQueues_43_reset = reset;
  assign taskQueues_43_io_connVec_0_push_valid = io_connPE_43_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_43_io_connVec_0_push_bits = io_connPE_43_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_43_io_connVec_0_pop_ready = io_connPE_43_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_43_io_connVec_1_push_valid = stealServers_43_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_43_io_connVec_1_push_bits = stealServers_43_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_43_io_connVec_1_pop_ready = stealServers_43_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_44_clock = clock;
  assign taskQueues_44_reset = reset;
  assign taskQueues_44_io_connVec_0_push_valid = io_connPE_44_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_44_io_connVec_0_push_bits = io_connPE_44_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_44_io_connVec_0_pop_ready = io_connPE_44_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_44_io_connVec_1_push_valid = stealServers_44_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_44_io_connVec_1_push_bits = stealServers_44_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_44_io_connVec_1_pop_ready = stealServers_44_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_45_clock = clock;
  assign taskQueues_45_reset = reset;
  assign taskQueues_45_io_connVec_0_push_valid = io_connPE_45_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_45_io_connVec_0_push_bits = io_connPE_45_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_45_io_connVec_0_pop_ready = io_connPE_45_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_45_io_connVec_1_push_valid = stealServers_45_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_45_io_connVec_1_push_bits = stealServers_45_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_45_io_connVec_1_pop_ready = stealServers_45_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_46_clock = clock;
  assign taskQueues_46_reset = reset;
  assign taskQueues_46_io_connVec_0_push_valid = io_connPE_46_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_46_io_connVec_0_push_bits = io_connPE_46_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_46_io_connVec_0_pop_ready = io_connPE_46_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_46_io_connVec_1_push_valid = stealServers_46_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_46_io_connVec_1_push_bits = stealServers_46_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_46_io_connVec_1_pop_ready = stealServers_46_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_47_clock = clock;
  assign taskQueues_47_reset = reset;
  assign taskQueues_47_io_connVec_0_push_valid = io_connPE_47_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_47_io_connVec_0_push_bits = io_connPE_47_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_47_io_connVec_0_pop_ready = io_connPE_47_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_47_io_connVec_1_push_valid = stealServers_47_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_47_io_connVec_1_push_bits = stealServers_47_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_47_io_connVec_1_pop_ready = stealServers_47_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_48_clock = clock;
  assign taskQueues_48_reset = reset;
  assign taskQueues_48_io_connVec_0_push_valid = io_connPE_48_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_48_io_connVec_0_push_bits = io_connPE_48_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_48_io_connVec_0_pop_ready = io_connPE_48_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_48_io_connVec_1_push_valid = stealServers_48_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_48_io_connVec_1_push_bits = stealServers_48_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_48_io_connVec_1_pop_ready = stealServers_48_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_49_clock = clock;
  assign taskQueues_49_reset = reset;
  assign taskQueues_49_io_connVec_0_push_valid = io_connPE_49_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_49_io_connVec_0_push_bits = io_connPE_49_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_49_io_connVec_0_pop_ready = io_connPE_49_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_49_io_connVec_1_push_valid = stealServers_49_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_49_io_connVec_1_push_bits = stealServers_49_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_49_io_connVec_1_pop_ready = stealServers_49_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_50_clock = clock;
  assign taskQueues_50_reset = reset;
  assign taskQueues_50_io_connVec_0_push_valid = io_connPE_50_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_50_io_connVec_0_push_bits = io_connPE_50_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_50_io_connVec_0_pop_ready = io_connPE_50_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_50_io_connVec_1_push_valid = stealServers_50_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_50_io_connVec_1_push_bits = stealServers_50_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_50_io_connVec_1_pop_ready = stealServers_50_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_51_clock = clock;
  assign taskQueues_51_reset = reset;
  assign taskQueues_51_io_connVec_0_push_valid = io_connPE_51_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_51_io_connVec_0_push_bits = io_connPE_51_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_51_io_connVec_0_pop_ready = io_connPE_51_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_51_io_connVec_1_push_valid = stealServers_51_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_51_io_connVec_1_push_bits = stealServers_51_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_51_io_connVec_1_pop_ready = stealServers_51_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_52_clock = clock;
  assign taskQueues_52_reset = reset;
  assign taskQueues_52_io_connVec_0_push_valid = io_connPE_52_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_52_io_connVec_0_push_bits = io_connPE_52_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_52_io_connVec_0_pop_ready = io_connPE_52_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_52_io_connVec_1_push_valid = stealServers_52_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_52_io_connVec_1_push_bits = stealServers_52_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_52_io_connVec_1_pop_ready = stealServers_52_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_53_clock = clock;
  assign taskQueues_53_reset = reset;
  assign taskQueues_53_io_connVec_0_push_valid = io_connPE_53_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_53_io_connVec_0_push_bits = io_connPE_53_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_53_io_connVec_0_pop_ready = io_connPE_53_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_53_io_connVec_1_push_valid = stealServers_53_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_53_io_connVec_1_push_bits = stealServers_53_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_53_io_connVec_1_pop_ready = stealServers_53_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_54_clock = clock;
  assign taskQueues_54_reset = reset;
  assign taskQueues_54_io_connVec_0_push_valid = io_connPE_54_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_54_io_connVec_0_push_bits = io_connPE_54_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_54_io_connVec_0_pop_ready = io_connPE_54_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_54_io_connVec_1_push_valid = stealServers_54_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_54_io_connVec_1_push_bits = stealServers_54_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_54_io_connVec_1_pop_ready = stealServers_54_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_55_clock = clock;
  assign taskQueues_55_reset = reset;
  assign taskQueues_55_io_connVec_0_push_valid = io_connPE_55_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_55_io_connVec_0_push_bits = io_connPE_55_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_55_io_connVec_0_pop_ready = io_connPE_55_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_55_io_connVec_1_push_valid = stealServers_55_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_55_io_connVec_1_push_bits = stealServers_55_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_55_io_connVec_1_pop_ready = stealServers_55_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_56_clock = clock;
  assign taskQueues_56_reset = reset;
  assign taskQueues_56_io_connVec_0_push_valid = io_connPE_56_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_56_io_connVec_0_push_bits = io_connPE_56_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_56_io_connVec_0_pop_ready = io_connPE_56_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_56_io_connVec_1_push_valid = stealServers_56_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_56_io_connVec_1_push_bits = stealServers_56_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_56_io_connVec_1_pop_ready = stealServers_56_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_57_clock = clock;
  assign taskQueues_57_reset = reset;
  assign taskQueues_57_io_connVec_0_push_valid = io_connPE_57_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_57_io_connVec_0_push_bits = io_connPE_57_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_57_io_connVec_0_pop_ready = io_connPE_57_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_57_io_connVec_1_push_valid = stealServers_57_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_57_io_connVec_1_push_bits = stealServers_57_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_57_io_connVec_1_pop_ready = stealServers_57_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_58_clock = clock;
  assign taskQueues_58_reset = reset;
  assign taskQueues_58_io_connVec_0_push_valid = io_connPE_58_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_58_io_connVec_0_push_bits = io_connPE_58_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_58_io_connVec_0_pop_ready = io_connPE_58_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_58_io_connVec_1_push_valid = stealServers_58_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_58_io_connVec_1_push_bits = stealServers_58_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_58_io_connVec_1_pop_ready = stealServers_58_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_59_clock = clock;
  assign taskQueues_59_reset = reset;
  assign taskQueues_59_io_connVec_0_push_valid = io_connPE_59_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_59_io_connVec_0_push_bits = io_connPE_59_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_59_io_connVec_0_pop_ready = io_connPE_59_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_59_io_connVec_1_push_valid = stealServers_59_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_59_io_connVec_1_push_bits = stealServers_59_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_59_io_connVec_1_pop_ready = stealServers_59_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_60_clock = clock;
  assign taskQueues_60_reset = reset;
  assign taskQueues_60_io_connVec_0_push_valid = io_connPE_60_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_60_io_connVec_0_push_bits = io_connPE_60_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_60_io_connVec_0_pop_ready = io_connPE_60_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_60_io_connVec_1_push_valid = stealServers_60_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_60_io_connVec_1_push_bits = stealServers_60_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_60_io_connVec_1_pop_ready = stealServers_60_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_61_clock = clock;
  assign taskQueues_61_reset = reset;
  assign taskQueues_61_io_connVec_0_push_valid = io_connPE_61_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_61_io_connVec_0_push_bits = io_connPE_61_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_61_io_connVec_0_pop_ready = io_connPE_61_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_61_io_connVec_1_push_valid = stealServers_61_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_61_io_connVec_1_push_bits = stealServers_61_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_61_io_connVec_1_pop_ready = stealServers_61_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_62_clock = clock;
  assign taskQueues_62_reset = reset;
  assign taskQueues_62_io_connVec_0_push_valid = io_connPE_62_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_62_io_connVec_0_push_bits = io_connPE_62_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_62_io_connVec_0_pop_ready = io_connPE_62_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_62_io_connVec_1_push_valid = stealServers_62_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_62_io_connVec_1_push_bits = stealServers_62_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_62_io_connVec_1_pop_ready = stealServers_62_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_63_clock = clock;
  assign taskQueues_63_reset = reset;
  assign taskQueues_63_io_connVec_0_push_valid = io_connPE_63_push_valid; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_63_io_connVec_0_push_bits = io_connPE_63_push_bits; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_63_io_connVec_0_pop_ready = io_connPE_63_pop_ready; // @[stealNW_TQ.scala 62:37]
  assign taskQueues_63_io_connVec_1_push_valid = stealServers_63_io_connQ_push_valid; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_63_io_connVec_1_push_bits = stealServers_63_io_connQ_push_bits; // @[stealNW_TQ.scala 69:37]
  assign taskQueues_63_io_connVec_1_pop_ready = stealServers_63_io_connQ_pop_ready; // @[stealNW_TQ.scala 69:37]
endmodule
module Queue(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [5:0] io_enq_bits_addr,
  input        io_deq_ready,
  output       io_deq_valid,
  output [5:0] io_deq_bits_addr
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [5:0] ram_addr [0:3]; // @[Decoupled.scala 275:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[Decoupled.scala 275:95]
  wire [1:0] ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 275:95]
  wire [5:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 275:95]
  wire [5:0] ram_addr_MPORT_data; // @[Decoupled.scala 275:95]
  wire [1:0] ram_addr_MPORT_addr; // @[Decoupled.scala 275:95]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 275:95]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 275:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 278:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 279:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 280:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 281:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 52:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 52:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 275:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = enq_ptr_value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 305:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 304:19]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 312:17]
  always @(posedge clock) begin
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 275:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 288:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 292:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 278:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 278:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 295:27]
      maybe_full <= do_enq; // @[Decoupled.scala 296:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[5:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_2(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_data,
  input  [7:0]  io_enq_bits_strb,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_data,
  output [7:0]  io_deq_bits_strb
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_data [0:3]; // @[Decoupled.scala 275:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[Decoupled.scala 275:95]
  wire [1:0] ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 275:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 275:95]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 275:95]
  wire [1:0] ram_data_MPORT_addr; // @[Decoupled.scala 275:95]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 275:95]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 275:95]
  reg [7:0] ram_strb [0:3]; // @[Decoupled.scala 275:95]
  wire  ram_strb_io_deq_bits_MPORT_en; // @[Decoupled.scala 275:95]
  wire [1:0] ram_strb_io_deq_bits_MPORT_addr; // @[Decoupled.scala 275:95]
  wire [7:0] ram_strb_io_deq_bits_MPORT_data; // @[Decoupled.scala 275:95]
  wire [7:0] ram_strb_MPORT_data; // @[Decoupled.scala 275:95]
  wire [1:0] ram_strb_MPORT_addr; // @[Decoupled.scala 275:95]
  wire  ram_strb_MPORT_mask; // @[Decoupled.scala 275:95]
  wire  ram_strb_MPORT_en; // @[Decoupled.scala 275:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 278:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 279:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 280:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 281:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 52:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 52:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 275:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_strb_io_deq_bits_MPORT_en = 1'h1;
  assign ram_strb_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_strb_io_deq_bits_MPORT_data = ram_strb[ram_strb_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 275:95]
  assign ram_strb_MPORT_data = io_enq_bits_strb;
  assign ram_strb_MPORT_addr = enq_ptr_value;
  assign ram_strb_MPORT_mask = 1'h1;
  assign ram_strb_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 305:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 304:19]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 312:17]
  assign io_deq_bits_strb = ram_strb_io_deq_bits_MPORT_data; // @[Decoupled.scala 312:17]
  always @(posedge clock) begin
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 275:95]
    end
    if (ram_strb_MPORT_en & ram_strb_MPORT_mask) begin
      ram_strb[ram_strb_MPORT_addr] <= ram_strb_MPORT_data; // @[Decoupled.scala 275:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 288:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 292:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 278:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 278:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 295:27]
      maybe_full <= do_enq; // @[Decoupled.scala 296:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_strb[initvar] = _RAND_1[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_3(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [255:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [255:0] io_deq_bits,
  output [4:0]   io_count
);
`ifdef RANDOMIZE_MEM_INIT
  reg [255:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [255:0] ram [0:15]; // @[Decoupled.scala 275:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 275:95]
  wire [3:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 275:95]
  wire [255:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 275:95]
  wire [255:0] ram_MPORT_data; // @[Decoupled.scala 275:95]
  wire [3:0] ram_MPORT_addr; // @[Decoupled.scala 275:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 275:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 275:95]
  reg [3:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [3:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 278:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 279:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 280:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 281:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 52:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 52:35]
  wire [3:0] _value_T_1 = enq_ptr_value + 4'h1; // @[Counter.scala 77:24]
  wire [3:0] _value_T_3 = deq_ptr_value + 4'h1; // @[Counter.scala 77:24]
  wire [3:0] ptr_diff = enq_ptr_value - deq_ptr_value; // @[Decoupled.scala 328:32]
  wire [4:0] _io_count_T_1 = maybe_full & ptr_match ? 5'h10 : 5'h0; // @[Decoupled.scala 331:20]
  wire [4:0] _GEN_11 = {{1'd0}, ptr_diff}; // @[Decoupled.scala 331:62]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 275:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 305:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 304:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 312:17]
  assign io_count = _io_count_T_1 | _GEN_11; // @[Decoupled.scala 331:62]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 275:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 4'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 288:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 4'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 292:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 278:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 278:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 295:27]
      maybe_full <= do_enq; // @[Decoupled.scala 296:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {8{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram[initvar] = _RAND_0[255:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module virtualStealServer(
  input          clock,
  input          reset,
  input          io_connNetwork_ctrl_serveStealReq_ready,
  output         io_connNetwork_ctrl_serveStealReq_valid,
  output         io_connNetwork_data_availableTask_ready,
  input          io_connNetwork_data_availableTask_valid,
  input  [255:0] io_connNetwork_data_availableTask_bits,
  input          io_connNetwork_data_qOutTask_ready,
  output         io_connNetwork_data_qOutTask_valid,
  output [255:0] io_connNetwork_data_qOutTask_bits,
  output         io_axi_mgmt_ARREADY,
  input          io_axi_mgmt_ARVALID,
  input  [5:0]   io_axi_mgmt_ARADDR,
  input          io_axi_mgmt_RREADY,
  output         io_axi_mgmt_RVALID,
  output [63:0]  io_axi_mgmt_RDATA,
  output         io_axi_mgmt_AWREADY,
  input          io_axi_mgmt_AWVALID,
  input  [5:0]   io_axi_mgmt_AWADDR,
  output         io_axi_mgmt_WREADY,
  input          io_axi_mgmt_WVALID,
  input  [63:0]  io_axi_mgmt_WDATA,
  input  [7:0]   io_axi_mgmt_WSTRB,
  input          io_axi_mgmt_BREADY,
  output         io_axi_mgmt_BVALID,
  input          io_read_address_ready,
  output         io_read_address_valid,
  output [63:0]  io_read_address_bits,
  output         io_read_data_ready,
  input          io_read_data_valid,
  input  [255:0] io_read_data_bits,
  output [3:0]   io_read_burst_len,
  input          io_write_address_ready,
  output         io_write_address_valid,
  output [63:0]  io_write_address_bits,
  input          io_write_data_ready,
  output         io_write_data_valid,
  output [255:0] io_write_data_bits,
  output [3:0]   io_write_burst_len,
  output         io_write_last,
  input          io_ntwDataUnitOccupancy
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  rdReq__deq_clock; // @[Decoupled.scala 377:21]
  wire  rdReq__deq_reset; // @[Decoupled.scala 377:21]
  wire  rdReq__deq_io_enq_ready; // @[Decoupled.scala 377:21]
  wire  rdReq__deq_io_enq_valid; // @[Decoupled.scala 377:21]
  wire [5:0] rdReq__deq_io_enq_bits_addr; // @[Decoupled.scala 377:21]
  wire  rdReq__deq_io_deq_ready; // @[Decoupled.scala 377:21]
  wire  rdReq__deq_io_deq_valid; // @[Decoupled.scala 377:21]
  wire [5:0] rdReq__deq_io_deq_bits_addr; // @[Decoupled.scala 377:21]
  wire  wrReq__deq_clock; // @[Decoupled.scala 377:21]
  wire  wrReq__deq_reset; // @[Decoupled.scala 377:21]
  wire  wrReq__deq_io_enq_ready; // @[Decoupled.scala 377:21]
  wire  wrReq__deq_io_enq_valid; // @[Decoupled.scala 377:21]
  wire [5:0] wrReq__deq_io_enq_bits_addr; // @[Decoupled.scala 377:21]
  wire  wrReq__deq_io_deq_ready; // @[Decoupled.scala 377:21]
  wire  wrReq__deq_io_deq_valid; // @[Decoupled.scala 377:21]
  wire [5:0] wrReq__deq_io_deq_bits_addr; // @[Decoupled.scala 377:21]
  wire  wrReqData__deq_clock; // @[Decoupled.scala 377:21]
  wire  wrReqData__deq_reset; // @[Decoupled.scala 377:21]
  wire  wrReqData__deq_io_enq_ready; // @[Decoupled.scala 377:21]
  wire  wrReqData__deq_io_enq_valid; // @[Decoupled.scala 377:21]
  wire [63:0] wrReqData__deq_io_enq_bits_data; // @[Decoupled.scala 377:21]
  wire [7:0] wrReqData__deq_io_enq_bits_strb; // @[Decoupled.scala 377:21]
  wire  wrReqData__deq_io_deq_ready; // @[Decoupled.scala 377:21]
  wire  wrReqData__deq_io_deq_valid; // @[Decoupled.scala 377:21]
  wire [63:0] wrReqData__deq_io_deq_bits_data; // @[Decoupled.scala 377:21]
  wire [7:0] wrReqData__deq_io_deq_bits_strb; // @[Decoupled.scala 377:21]
  wire  taskQueueBuffer_clock; // @[virtualStealServer.scala 81:43]
  wire  taskQueueBuffer_reset; // @[virtualStealServer.scala 81:43]
  wire  taskQueueBuffer_io_enq_ready; // @[virtualStealServer.scala 81:43]
  wire  taskQueueBuffer_io_enq_valid; // @[virtualStealServer.scala 81:43]
  wire [255:0] taskQueueBuffer_io_enq_bits; // @[virtualStealServer.scala 81:43]
  wire  taskQueueBuffer_io_deq_ready; // @[virtualStealServer.scala 81:43]
  wire  taskQueueBuffer_io_deq_valid; // @[virtualStealServer.scala 81:43]
  wire [255:0] taskQueueBuffer_io_deq_bits; // @[virtualStealServer.scala 81:43]
  wire [4:0] taskQueueBuffer_io_count; // @[virtualStealServer.scala 81:43]
  wire  rdReq__valid = rdReq__deq_io_deq_valid; // @[Decoupled.scala 417:19 419:15]
  wire  rdReq = rdReq__valid & io_axi_mgmt_RREADY; // @[RegisterBlock.scala 210:44]
  wire [5:0] rdReq__bits_addr = rdReq__deq_io_deq_bits_addr; // @[Decoupled.scala 417:19 418:14]
  wire [5:0] rdAddr = rdReq__bits_addr & 6'h38; // @[RegisterBlock.scala 214:48]
  wire  wrReq__valid = wrReq__deq_io_deq_valid; // @[Decoupled.scala 417:19 419:15]
  wire  wrReqData__valid = wrReqData__deq_io_deq_valid; // @[Decoupled.scala 417:19 419:15]
  wire  wrReq = wrReq__valid & wrReqData__valid & io_axi_mgmt_BREADY; // @[RegisterBlock.scala 241:63]
  wire [5:0] wrReq__bits_addr = wrReq__deq_io_deq_bits_addr; // @[Decoupled.scala 417:19 418:14]
  wire [5:0] wrAddr = wrReq__bits_addr & 6'h38; // @[RegisterBlock.scala 243:48]
  reg [63:0] rAddr; // @[virtualStealServer.scala 65:44]
  reg [63:0] rPause; // @[virtualStealServer.scala 66:44]
  reg [63:0] procInterrupt; // @[virtualStealServer.scala 67:44]
  reg [63:0] maxLength; // @[virtualStealServer.scala 68:44]
  reg [3:0] stateReg; // @[virtualStealServer.scala 69:44]
  reg [63:0] contentionCounter; // @[virtualStealServer.scala 71:44]
  reg  networkCongested; // @[virtualStealServer.scala 73:44]
  reg [63:0] fifoTailReg; // @[virtualStealServer.scala 77:44]
  reg [63:0] fifoHeadReg; // @[virtualStealServer.scala 78:44]
  reg  popOrPush; // @[virtualStealServer.scala 79:44]
  reg [4:0] memDataCounter; // @[virtualStealServer.scala 82:44]
  wire [63:0] _contentionCounter_T_1 = contentionCounter + 64'h1; // @[virtualStealServer.scala 98:52]
  wire  _T_2 = contentionCounter != 64'h0; // @[virtualStealServer.scala 99:38]
  wire [63:0] _contentionCounter_T_3 = contentionCounter - 64'h1; // @[virtualStealServer.scala 101:52]
  wire [63:0] _T_9 = 64'h37 - 64'h0; // @[virtualStealServer.scala 122:54]
  wire  _GEN_2 = contentionCounter < _T_9 ? 1'h0 : networkCongested; // @[virtualStealServer.scala 122:63 123:26 125:26]
  wire  _GEN_3 = contentionCounter >= 64'h37 | _GEN_2; // @[virtualStealServer.scala 120:58 121:26]
  wire [63:0] _currLen_T_1 = fifoTailReg - fifoHeadReg; // @[virtualStealServer.scala 359:32]
  wire [63:0] _currLen_T_3 = maxLength - fifoHeadReg; // @[virtualStealServer.scala 364:30]
  wire [63:0] _currLen_T_5 = _currLen_T_3 + fifoTailReg; // @[virtualStealServer.scala 364:44]
  reg [63:0] lengthHistroy; // @[virtualStealServer.scala 355:32]
  wire [63:0] _currLen_T_7 = lengthHistroy + 64'h1; // @[virtualStealServer.scala 377:38]
  wire [63:0] _GEN_138 = popOrPush ? 64'h0 : _currLen_T_7; // @[virtualStealServer.scala 371:24 373:21 377:21]
  wire [63:0] _GEN_139 = fifoTailReg < fifoHeadReg ? _currLen_T_5 : _GEN_138; // @[virtualStealServer.scala 362:42 364:17]
  wire [63:0] currLen = fifoTailReg > fifoHeadReg ? _currLen_T_1 : _GEN_139; // @[virtualStealServer.scala 357:36 359:17]
  wire [63:0] _T_15 = 64'h10 + currLen; // @[virtualStealServer.scala 132:79]
  wire  _T_20 = ~networkCongested; // @[virtualStealServer.scala 145:20]
  wire [3:0] _GEN_4 = procInterrupt != 64'h0 ? 4'ha : stateReg; // @[virtualStealServer.scala 153:42 155:22 69:44]
  wire [63:0] _GEN_5 = procInterrupt != 64'h0 ? 64'hffffffffffffffff : rPause; // @[virtualStealServer.scala 153:42 156:22 66:44]
  wire [3:0] _GEN_6 = _T_20 & taskQueueBuffer_io_count != 5'h0 ? 4'h7 : _GEN_4; // @[virtualStealServer.scala 149:74 151:22]
  wire [63:0] _GEN_7 = _T_20 & taskQueueBuffer_io_count != 5'h0 ? rPause : _GEN_5; // @[virtualStealServer.scala 149:74 66:44]
  wire [3:0] _GEN_8 = ~networkCongested & currLen != 64'h0 & taskQueueBuffer_io_count == 5'h0 ? 4'h6 : _GEN_6; // @[virtualStealServer.scala 145:93 147:22]
  wire [63:0] _GEN_9 = ~networkCongested & currLen != 64'h0 & taskQueueBuffer_io_count == 5'h0 ? rPause : _GEN_7; // @[virtualStealServer.scala 145:93 66:44]
  wire [3:0] _GEN_10 = networkCongested ? 4'h2 : _GEN_8; // @[virtualStealServer.scala 141:37 143:22]
  wire [63:0] _GEN_11 = networkCongested ? rPause : _GEN_9; // @[virtualStealServer.scala 141:37 66:44]
  wire [63:0] _GEN_13 = networkCongested & taskQueueBuffer_io_count == 5'h10 ? rPause : _GEN_11; // @[virtualStealServer.scala 137:74 66:44]
  wire [63:0] _GEN_15 = currLen == maxLength & networkCongested | maxLength < _T_15 ? 64'hffffffffffffffff : _GEN_13; // @[virtualStealServer.scala 132:90 135:22]
  wire  _T_29 = stateReg == 4'h2; // @[virtualStealServer.scala 160:25]
  wire [3:0] _GEN_16 = _T_20 ? 4'h0 : stateReg; // @[virtualStealServer.scala 170:38 172:22 69:44]
  wire [3:0] _GEN_17 = io_connNetwork_data_availableTask_valid & networkCongested ? 4'h2 : _GEN_16; // @[virtualStealServer.scala 166:80 168:22]
  wire  _T_34 = stateReg == 4'h4; // @[virtualStealServer.scala 176:25]
  wire [3:0] _GEN_19 = io_write_address_ready ? 4'h3 : stateReg; // @[virtualStealServer.scala 178:37 179:22 69:44]
  wire [4:0] _GEN_20 = io_write_address_ready ? 5'h10 : memDataCounter; // @[virtualStealServer.scala 178:37 180:28 82:44]
  wire  _T_35 = stateReg == 4'h3; // @[virtualStealServer.scala 183:25]
  wire  _T_36 = memDataCounter == 5'h1; // @[virtualStealServer.scala 185:52]
  wire [63:0] _T_39 = maxLength - 64'h1; // @[virtualStealServer.scala 189:42]
  wire [63:0] _fifoTailReg_T_1 = fifoTailReg + 64'h1; // @[virtualStealServer.scala 190:44]
  wire [63:0] _GEN_21 = fifoTailReg < _T_39 ? _fifoTailReg_T_1 : 64'h0; // @[virtualStealServer.scala 189:48 190:29 192:29]
  wire [4:0] _memDataCounter_T_1 = memDataCounter - 5'h1; // @[virtualStealServer.scala 196:46]
  wire [4:0] _GEN_23 = io_write_data_ready ? _memDataCounter_T_1 : memDataCounter; // @[virtualStealServer.scala 195:40 196:28 82:44]
  wire [63:0] _GEN_24 = io_write_data_ready ? _GEN_21 : fifoTailReg; // @[virtualStealServer.scala 195:40 77:44]
  wire [3:0] _GEN_25 = io_write_data_ready & memDataCounter == 5'h1 ? 4'h0 : stateReg; // @[virtualStealServer.scala 185:60 186:22 69:44]
  wire  _GEN_26 = io_write_data_ready & memDataCounter == 5'h1 ? 1'h0 : popOrPush; // @[virtualStealServer.scala 185:60 187:23 79:44]
  wire [63:0] _GEN_27 = io_write_data_ready & memDataCounter == 5'h1 ? _GEN_21 : _GEN_24; // @[virtualStealServer.scala 185:60]
  wire [4:0] _GEN_28 = io_write_data_ready & memDataCounter == 5'h1 ? memDataCounter : _GEN_23; // @[virtualStealServer.scala 185:60 82:44]
  wire  _T_44 = stateReg == 4'h6; // @[virtualStealServer.scala 204:25]
  wire  _memDataCounter_T_2 = currLen < 64'h10; // @[virtualStealServer.scala 208:43]
  wire [63:0] _memDataCounter_T_3 = currLen < 64'h10 ? currLen : 64'h10; // @[virtualStealServer.scala 208:34]
  wire [3:0] _GEN_29 = io_read_address_ready ? 4'h5 : stateReg; // @[virtualStealServer.scala 206:36 207:22 69:44]
  wire [63:0] _GEN_30 = io_read_address_ready ? _memDataCounter_T_3 : {{59'd0}, memDataCounter}; // @[virtualStealServer.scala 206:36 208:28 82:44]
  wire  _T_45 = stateReg == 4'h5; // @[virtualStealServer.scala 211:25]
  wire [63:0] _fifoHeadReg_T_1 = fifoHeadReg + 64'h1; // @[virtualStealServer.scala 218:44]
  wire [63:0] _GEN_31 = fifoHeadReg < _T_39 ? _fifoHeadReg_T_1 : 64'h0; // @[virtualStealServer.scala 217:48 218:29 220:29]
  wire [4:0] _GEN_33 = io_read_data_valid ? _memDataCounter_T_1 : memDataCounter; // @[virtualStealServer.scala 222:39 223:28 82:44]
  wire [63:0] _GEN_34 = io_read_data_valid ? _GEN_31 : fifoHeadReg; // @[virtualStealServer.scala 222:39 78:44]
  wire [3:0] _GEN_35 = io_read_data_valid & _T_36 ? 4'h8 : stateReg; // @[virtualStealServer.scala 213:59 214:22 69:44]
  wire  _GEN_36 = io_read_data_valid & _T_36 | popOrPush; // @[virtualStealServer.scala 213:59 215:23 79:44]
  wire [63:0] _GEN_37 = io_read_data_valid & _T_36 ? _GEN_31 : _GEN_34; // @[virtualStealServer.scala 213:59]
  wire [4:0] _GEN_38 = io_read_data_valid & _T_36 ? memDataCounter : _GEN_33; // @[virtualStealServer.scala 213:59 82:44]
  wire  _T_54 = stateReg == 4'h7; // @[virtualStealServer.scala 231:25]
  wire [2:0] _GEN_39 = networkCongested ? 3'h0 : 3'h7; // @[virtualStealServer.scala 235:37 236:22 238:22]
  wire [2:0] _GEN_40 = io_connNetwork_data_qOutTask_ready ? 3'h0 : _GEN_39; // @[virtualStealServer.scala 233:49 234:22]
  wire  _T_55 = stateReg == 4'h8; // @[virtualStealServer.scala 241:25]
  wire [3:0] _GEN_41 = networkCongested ? 4'h0 : stateReg; // @[virtualStealServer.scala 247:37 249:22 69:44]
  wire [3:0] _GEN_42 = io_connNetwork_ctrl_serveStealReq_ready ? 4'h7 : _GEN_41; // @[virtualStealServer.scala 243:54 245:22]
  wire  _T_57 = rPause == 64'h0; // @[virtualStealServer.scala 255:21]
  wire [3:0] _GEN_43 = rPause == 64'h0 ? 4'h0 : 4'h9; // @[virtualStealServer.scala 255:33 257:22 261:22]
  wire [3:0] _GEN_44 = _T_57 ? 4'h0 : 4'ha; // @[virtualStealServer.scala 267:33 268:22 270:22]
  wire [3:0] _GEN_45 = stateReg == 4'ha ? _GEN_44 : stateReg; // @[virtualStealServer.scala 265:57 69:44]
  wire [3:0] _GEN_46 = stateReg == 4'h9 ? _GEN_43 : _GEN_45; // @[virtualStealServer.scala 253:46]
  wire [3:0] _GEN_47 = stateReg == 4'h8 ? _GEN_42 : _GEN_46; // @[virtualStealServer.scala 241:54]
  wire [3:0] _GEN_48 = stateReg == 4'h7 ? {{1'd0}, _GEN_40} : _GEN_47; // @[virtualStealServer.scala 231:48]
  wire [3:0] _GEN_49 = stateReg == 4'h5 ? _GEN_35 : _GEN_48; // @[virtualStealServer.scala 211:46]
  wire  _GEN_50 = stateReg == 4'h5 ? _GEN_36 : popOrPush; // @[virtualStealServer.scala 211:46 79:44]
  wire [63:0] _GEN_51 = stateReg == 4'h5 ? _GEN_37 : fifoHeadReg; // @[virtualStealServer.scala 211:46 78:44]
  wire [4:0] _GEN_52 = stateReg == 4'h5 ? _GEN_38 : memDataCounter; // @[virtualStealServer.scala 211:46 82:44]
  wire [3:0] _GEN_53 = stateReg == 4'h6 ? _GEN_29 : _GEN_49; // @[virtualStealServer.scala 204:53]
  wire [63:0] _GEN_54 = stateReg == 4'h6 ? _GEN_30 : {{59'd0}, _GEN_52}; // @[virtualStealServer.scala 204:53]
  wire  _GEN_55 = stateReg == 4'h6 ? popOrPush : _GEN_50; // @[virtualStealServer.scala 204:53 79:44]
  wire [63:0] _GEN_56 = stateReg == 4'h6 ? fifoHeadReg : _GEN_51; // @[virtualStealServer.scala 204:53 78:44]
  wire [3:0] _GEN_57 = stateReg == 4'h3 ? _GEN_25 : _GEN_53; // @[virtualStealServer.scala 183:47]
  wire  _GEN_58 = stateReg == 4'h3 ? _GEN_26 : _GEN_55; // @[virtualStealServer.scala 183:47]
  wire [63:0] _GEN_59 = stateReg == 4'h3 ? _GEN_27 : fifoTailReg; // @[virtualStealServer.scala 183:47 77:44]
  wire [63:0] _GEN_60 = stateReg == 4'h3 ? {{59'd0}, _GEN_28} : _GEN_54; // @[virtualStealServer.scala 183:47]
  wire [63:0] _GEN_61 = stateReg == 4'h3 ? fifoHeadReg : _GEN_56; // @[virtualStealServer.scala 183:47 78:44]
  wire [63:0] _GEN_63 = stateReg == 4'h4 ? {{59'd0}, _GEN_20} : _GEN_60; // @[virtualStealServer.scala 176:54]
  wire  _GEN_64 = stateReg == 4'h4 ? popOrPush : _GEN_58; // @[virtualStealServer.scala 176:54 79:44]
  wire [63:0] _GEN_65 = stateReg == 4'h4 ? fifoTailReg : _GEN_59; // @[virtualStealServer.scala 176:54 77:44]
  wire [63:0] _GEN_66 = stateReg == 4'h4 ? fifoHeadReg : _GEN_61; // @[virtualStealServer.scala 176:54 78:44]
  wire [63:0] _GEN_68 = stateReg == 4'h2 ? {{59'd0}, memDataCounter} : _GEN_63; // @[virtualStealServer.scala 160:46 82:44]
  wire  _GEN_69 = stateReg == 4'h2 ? popOrPush : _GEN_64; // @[virtualStealServer.scala 160:46 79:44]
  wire [63:0] _GEN_70 = stateReg == 4'h2 ? fifoTailReg : _GEN_65; // @[virtualStealServer.scala 160:46 77:44]
  wire [63:0] _GEN_71 = stateReg == 4'h2 ? fifoHeadReg : _GEN_66; // @[virtualStealServer.scala 160:46 78:44]
  wire [63:0] _GEN_73 = stateReg == 4'h0 ? _GEN_15 : rPause; // @[virtualStealServer.scala 130:34 66:44]
  wire [63:0] _GEN_74 = stateReg == 4'h0 ? {{59'd0}, memDataCounter} : _GEN_68; // @[virtualStealServer.scala 130:34 82:44]
  wire  _GEN_75 = stateReg == 4'h0 ? popOrPush : _GEN_69; // @[virtualStealServer.scala 130:34 79:44]
  wire [63:0] _GEN_76 = stateReg == 4'h0 ? fifoTailReg : _GEN_70; // @[virtualStealServer.scala 130:34 77:44]
  wire [63:0] _GEN_77 = stateReg == 4'h0 ? fifoHeadReg : _GEN_71; // @[virtualStealServer.scala 130:34 78:44]
  wire [68:0] _GEN_166 = {fifoTailReg, 5'h0}; // @[virtualStealServer.scala 318:65]
  wire [70:0] _io_write_address_bits_T = {{2'd0}, _GEN_166}; // @[virtualStealServer.scala 318:65]
  wire [70:0] _GEN_167 = {{7'd0}, rAddr}; // @[virtualStealServer.scala 318:79]
  wire [70:0] _io_write_address_bits_T_2 = _io_write_address_bits_T + _GEN_167; // @[virtualStealServer.scala 318:79]
  wire [68:0] _GEN_168 = {fifoHeadReg, 5'h0}; // @[virtualStealServer.scala 333:65]
  wire [70:0] _io_read_address_bits_T = {{2'd0}, _GEN_168}; // @[virtualStealServer.scala 333:65]
  wire [70:0] _io_read_address_bits_T_2 = _io_read_address_bits_T + _GEN_167; // @[virtualStealServer.scala 333:79]
  wire [63:0] _io_read_burst_len_T_2 = currLen - 64'h1; // @[virtualStealServer.scala 334:79]
  wire [63:0] _io_read_burst_len_T_3 = _memDataCounter_T_2 ? _io_read_burst_len_T_2 : 64'hf; // @[virtualStealServer.scala 334:55]
  wire  _GEN_81 = _T_54 & io_connNetwork_data_qOutTask_ready; // @[virtualStealServer.scala 299:45 342:48 345:49]
  wire  _GEN_82 = _T_54 ? 1'h0 : _T_55; // @[virtualStealServer.scala 293:45 342:48]
  wire [255:0] _GEN_84 = _T_45 ? io_read_data_bits : 256'h0; // @[virtualStealServer.scala 297:45 336:46 339:49]
  wire  _GEN_85 = _T_45 & io_read_data_valid; // @[virtualStealServer.scala 296:45 336:46 340:49]
  wire  _GEN_86 = _T_45 ? 1'h0 : _T_54; // @[virtualStealServer.scala 289:45 336:46]
  wire  _GEN_87 = _T_45 ? 1'h0 : _GEN_81; // @[virtualStealServer.scala 299:45 336:46]
  wire  _GEN_88 = _T_45 ? 1'h0 : _GEN_82; // @[virtualStealServer.scala 293:45 336:46]
  wire [70:0] _GEN_90 = _T_44 ? _io_read_address_bits_T_2 : 71'h0; // @[virtualStealServer.scala 281:45 330:53 333:49]
  wire [63:0] _GEN_91 = _T_44 ? _io_read_burst_len_T_3 : 64'h0; // @[virtualStealServer.scala 304:45 330:53 334:49]
  wire  _GEN_92 = _T_44 ? 1'h0 : _T_45; // @[virtualStealServer.scala 282:45 330:53]
  wire [255:0] _GEN_93 = _T_44 ? 256'h0 : _GEN_84; // @[virtualStealServer.scala 297:45 330:53]
  wire  _GEN_94 = _T_44 ? 1'h0 : _GEN_85; // @[virtualStealServer.scala 296:45 330:53]
  wire  _GEN_95 = _T_44 ? 1'h0 : _GEN_86; // @[virtualStealServer.scala 289:45 330:53]
  wire  _GEN_96 = _T_44 ? 1'h0 : _GEN_87; // @[virtualStealServer.scala 299:45 330:53]
  wire  _GEN_97 = _T_44 ? 1'h0 : _GEN_88; // @[virtualStealServer.scala 293:45 330:53]
  wire  _GEN_99 = _T_35 ? io_write_data_ready : _GEN_96; // @[virtualStealServer.scala 321:47 324:49]
  wire  _GEN_100 = _T_35 & _T_36; // @[virtualStealServer.scala 303:45 321:47]
  wire  _GEN_101 = _T_35 ? 1'h0 : _T_44; // @[virtualStealServer.scala 280:45 321:47]
  wire [70:0] _GEN_102 = _T_35 ? 71'h0 : _GEN_90; // @[virtualStealServer.scala 281:45 321:47]
  wire [63:0] _GEN_103 = _T_35 ? 64'h0 : _GEN_91; // @[virtualStealServer.scala 304:45 321:47]
  wire  _GEN_104 = _T_35 ? 1'h0 : _GEN_92; // @[virtualStealServer.scala 282:45 321:47]
  wire [255:0] _GEN_105 = _T_35 ? 256'h0 : _GEN_93; // @[virtualStealServer.scala 297:45 321:47]
  wire  _GEN_106 = _T_35 ? 1'h0 : _GEN_94; // @[virtualStealServer.scala 296:45 321:47]
  wire  _GEN_107 = _T_35 ? 1'h0 : _GEN_95; // @[virtualStealServer.scala 289:45 321:47]
  wire  _GEN_108 = _T_35 ? 1'h0 : _GEN_97; // @[virtualStealServer.scala 293:45 321:47]
  wire [70:0] _GEN_110 = _T_34 ? _io_write_address_bits_T_2 : 71'h0; // @[virtualStealServer.scala 284:45 315:54 318:49]
  wire [3:0] _GEN_111 = _T_34 ? 4'hf : 4'h0; // @[virtualStealServer.scala 302:45 315:54 319:49]
  wire  _GEN_112 = _T_34 ? 1'h0 : _T_35; // @[virtualStealServer.scala 285:45 315:54]
  wire  _GEN_113 = _T_34 ? 1'h0 : _GEN_99; // @[virtualStealServer.scala 299:45 315:54]
  wire  _GEN_114 = _T_34 ? 1'h0 : _GEN_100; // @[virtualStealServer.scala 303:45 315:54]
  wire  _GEN_115 = _T_34 ? 1'h0 : _GEN_101; // @[virtualStealServer.scala 280:45 315:54]
  wire [70:0] _GEN_116 = _T_34 ? 71'h0 : _GEN_102; // @[virtualStealServer.scala 281:45 315:54]
  wire [63:0] _GEN_117 = _T_34 ? 64'h0 : _GEN_103; // @[virtualStealServer.scala 304:45 315:54]
  wire  _GEN_118 = _T_34 ? 1'h0 : _GEN_104; // @[virtualStealServer.scala 282:45 315:54]
  wire [255:0] _GEN_119 = _T_34 ? 256'h0 : _GEN_105; // @[virtualStealServer.scala 297:45 315:54]
  wire  _GEN_120 = _T_34 ? 1'h0 : _GEN_106; // @[virtualStealServer.scala 296:45 315:54]
  wire  _GEN_121 = _T_34 ? 1'h0 : _GEN_107; // @[virtualStealServer.scala 289:45 315:54]
  wire  _GEN_122 = _T_34 ? 1'h0 : _GEN_108; // @[virtualStealServer.scala 293:45 315:54]
  wire [70:0] _GEN_127 = _T_29 ? 71'h0 : _GEN_110; // @[virtualStealServer.scala 309:40 284:45]
  wire [70:0] _GEN_133 = _T_29 ? 71'h0 : _GEN_116; // @[virtualStealServer.scala 309:40 281:45]
  wire [63:0] _GEN_134 = _T_29 ? 64'h0 : _GEN_117; // @[virtualStealServer.scala 309:40 304:45]
  wire [63:0] _GEN_143 = 6'h0 == rdAddr ? rPause : 64'hffffffffffffffff; // @[RegisterBlock.scala 220:10 224:38 225:16]
  wire [63:0] _GEN_144 = 6'h8 == rdAddr ? rAddr : _GEN_143; // @[RegisterBlock.scala 224:38 225:16]
  wire [63:0] _GEN_145 = 6'h10 == rdAddr ? maxLength : _GEN_144; // @[RegisterBlock.scala 224:38 225:16]
  wire [63:0] _GEN_146 = 6'h18 == rdAddr ? fifoTailReg : _GEN_145; // @[RegisterBlock.scala 224:38 225:16]
  wire [63:0] _GEN_147 = 6'h20 == rdAddr ? fifoHeadReg : _GEN_146; // @[RegisterBlock.scala 224:38 225:16]
  wire  _T_77 = ~reset; // @[RegisterBlock.scala 182:11]
  wire [7:0] wrReqData__bits_strb = wrReqData__deq_io_deq_bits_strb; // @[Decoupled.scala 417:19 418:14]
  wire [63:0] wrReqData__bits_data = wrReqData__deq_io_deq_bits_data; // @[Decoupled.scala 417:19 418:14]
  wire [7:0] rPause_byte_wdata = wrReqData__bits_data[7:0]; // @[Interface.scala 257:33]
  wire [7:0] rPause_byte_original = rPause[7:0]; // @[Interface.scala 258:39]
  wire [7:0] _rPause_T_8 = wrReqData__bits_strb[0] ? rPause_byte_wdata : rPause_byte_original; // @[Interface.scala 259:14]
  wire [7:0] rPause_byte_wdata_1 = wrReqData__bits_data[15:8]; // @[Interface.scala 257:33]
  wire [7:0] rPause_byte_original_1 = rPause[15:8]; // @[Interface.scala 258:39]
  wire [7:0] _rPause_T_9 = wrReqData__bits_strb[1] ? rPause_byte_wdata_1 : rPause_byte_original_1; // @[Interface.scala 259:14]
  wire [7:0] rPause_byte_wdata_2 = wrReqData__bits_data[23:16]; // @[Interface.scala 257:33]
  wire [7:0] rPause_byte_original_2 = rPause[23:16]; // @[Interface.scala 258:39]
  wire [7:0] _rPause_T_10 = wrReqData__bits_strb[2] ? rPause_byte_wdata_2 : rPause_byte_original_2; // @[Interface.scala 259:14]
  wire [7:0] rPause_byte_wdata_3 = wrReqData__bits_data[31:24]; // @[Interface.scala 257:33]
  wire [7:0] rPause_byte_original_3 = rPause[31:24]; // @[Interface.scala 258:39]
  wire [7:0] _rPause_T_11 = wrReqData__bits_strb[3] ? rPause_byte_wdata_3 : rPause_byte_original_3; // @[Interface.scala 259:14]
  wire [7:0] rPause_byte_wdata_4 = wrReqData__bits_data[39:32]; // @[Interface.scala 257:33]
  wire [7:0] rPause_byte_original_4 = rPause[39:32]; // @[Interface.scala 258:39]
  wire [7:0] _rPause_T_12 = wrReqData__bits_strb[4] ? rPause_byte_wdata_4 : rPause_byte_original_4; // @[Interface.scala 259:14]
  wire [7:0] rPause_byte_wdata_5 = wrReqData__bits_data[47:40]; // @[Interface.scala 257:33]
  wire [7:0] rPause_byte_original_5 = rPause[47:40]; // @[Interface.scala 258:39]
  wire [7:0] _rPause_T_13 = wrReqData__bits_strb[5] ? rPause_byte_wdata_5 : rPause_byte_original_5; // @[Interface.scala 259:14]
  wire [7:0] rPause_byte_wdata_6 = wrReqData__bits_data[55:48]; // @[Interface.scala 257:33]
  wire [7:0] rPause_byte_original_6 = rPause[55:48]; // @[Interface.scala 258:39]
  wire [7:0] _rPause_T_14 = wrReqData__bits_strb[6] ? rPause_byte_wdata_6 : rPause_byte_original_6; // @[Interface.scala 259:14]
  wire [7:0] rPause_byte_wdata_7 = wrReqData__bits_data[63:56]; // @[Interface.scala 257:33]
  wire [7:0] rPause_byte_original_7 = rPause[63:56]; // @[Interface.scala 258:39]
  wire [7:0] _rPause_T_15 = wrReqData__bits_strb[7] ? rPause_byte_wdata_7 : rPause_byte_original_7; // @[Interface.scala 259:14]
  wire [63:0] _rPause_T_16 = {_rPause_T_15,_rPause_T_14,_rPause_T_13,_rPause_T_12,_rPause_T_11,_rPause_T_10,_rPause_T_9,
    _rPause_T_8}; // @[Interface.scala 262:7]
  wire [7:0] rAddr_byte_original = rAddr[7:0]; // @[Interface.scala 258:39]
  wire [7:0] _rAddr_T_8 = wrReqData__bits_strb[0] ? rPause_byte_wdata : rAddr_byte_original; // @[Interface.scala 259:14]
  wire [7:0] rAddr_byte_original_1 = rAddr[15:8]; // @[Interface.scala 258:39]
  wire [7:0] _rAddr_T_9 = wrReqData__bits_strb[1] ? rPause_byte_wdata_1 : rAddr_byte_original_1; // @[Interface.scala 259:14]
  wire [7:0] rAddr_byte_original_2 = rAddr[23:16]; // @[Interface.scala 258:39]
  wire [7:0] _rAddr_T_10 = wrReqData__bits_strb[2] ? rPause_byte_wdata_2 : rAddr_byte_original_2; // @[Interface.scala 259:14]
  wire [7:0] rAddr_byte_original_3 = rAddr[31:24]; // @[Interface.scala 258:39]
  wire [7:0] _rAddr_T_11 = wrReqData__bits_strb[3] ? rPause_byte_wdata_3 : rAddr_byte_original_3; // @[Interface.scala 259:14]
  wire [7:0] rAddr_byte_original_4 = rAddr[39:32]; // @[Interface.scala 258:39]
  wire [7:0] _rAddr_T_12 = wrReqData__bits_strb[4] ? rPause_byte_wdata_4 : rAddr_byte_original_4; // @[Interface.scala 259:14]
  wire [7:0] rAddr_byte_original_5 = rAddr[47:40]; // @[Interface.scala 258:39]
  wire [7:0] _rAddr_T_13 = wrReqData__bits_strb[5] ? rPause_byte_wdata_5 : rAddr_byte_original_5; // @[Interface.scala 259:14]
  wire [7:0] rAddr_byte_original_6 = rAddr[55:48]; // @[Interface.scala 258:39]
  wire [7:0] _rAddr_T_14 = wrReqData__bits_strb[6] ? rPause_byte_wdata_6 : rAddr_byte_original_6; // @[Interface.scala 259:14]
  wire [7:0] rAddr_byte_original_7 = rAddr[63:56]; // @[Interface.scala 258:39]
  wire [7:0] _rAddr_T_15 = wrReqData__bits_strb[7] ? rPause_byte_wdata_7 : rAddr_byte_original_7; // @[Interface.scala 259:14]
  wire [63:0] _rAddr_T_16 = {_rAddr_T_15,_rAddr_T_14,_rAddr_T_13,_rAddr_T_12,_rAddr_T_11,_rAddr_T_10,_rAddr_T_9,
    _rAddr_T_8}; // @[Interface.scala 262:7]
  wire [7:0] maxLength_byte_original = maxLength[7:0]; // @[Interface.scala 258:39]
  wire [7:0] _maxLength_T_8 = wrReqData__bits_strb[0] ? rPause_byte_wdata : maxLength_byte_original; // @[Interface.scala 259:14]
  wire [7:0] maxLength_byte_original_1 = maxLength[15:8]; // @[Interface.scala 258:39]
  wire [7:0] _maxLength_T_9 = wrReqData__bits_strb[1] ? rPause_byte_wdata_1 : maxLength_byte_original_1; // @[Interface.scala 259:14]
  wire [7:0] maxLength_byte_original_2 = maxLength[23:16]; // @[Interface.scala 258:39]
  wire [7:0] _maxLength_T_10 = wrReqData__bits_strb[2] ? rPause_byte_wdata_2 : maxLength_byte_original_2; // @[Interface.scala 259:14]
  wire [7:0] maxLength_byte_original_3 = maxLength[31:24]; // @[Interface.scala 258:39]
  wire [7:0] _maxLength_T_11 = wrReqData__bits_strb[3] ? rPause_byte_wdata_3 : maxLength_byte_original_3; // @[Interface.scala 259:14]
  wire [7:0] maxLength_byte_original_4 = maxLength[39:32]; // @[Interface.scala 258:39]
  wire [7:0] _maxLength_T_12 = wrReqData__bits_strb[4] ? rPause_byte_wdata_4 : maxLength_byte_original_4; // @[Interface.scala 259:14]
  wire [7:0] maxLength_byte_original_5 = maxLength[47:40]; // @[Interface.scala 258:39]
  wire [7:0] _maxLength_T_13 = wrReqData__bits_strb[5] ? rPause_byte_wdata_5 : maxLength_byte_original_5; // @[Interface.scala 259:14]
  wire [7:0] maxLength_byte_original_6 = maxLength[55:48]; // @[Interface.scala 258:39]
  wire [7:0] _maxLength_T_14 = wrReqData__bits_strb[6] ? rPause_byte_wdata_6 : maxLength_byte_original_6; // @[Interface.scala 259:14]
  wire [7:0] maxLength_byte_original_7 = maxLength[63:56]; // @[Interface.scala 258:39]
  wire [7:0] _maxLength_T_15 = wrReqData__bits_strb[7] ? rPause_byte_wdata_7 : maxLength_byte_original_7; // @[Interface.scala 259:14]
  wire [63:0] _maxLength_T_16 = {_maxLength_T_15,_maxLength_T_14,_maxLength_T_13,_maxLength_T_12,_maxLength_T_11,
    _maxLength_T_10,_maxLength_T_9,_maxLength_T_8}; // @[Interface.scala 262:7]
  wire [7:0] fifoTailReg_byte_original = fifoTailReg[7:0]; // @[Interface.scala 258:39]
  wire [7:0] _fifoTailReg_T_12 = wrReqData__bits_strb[0] ? rPause_byte_wdata : fifoTailReg_byte_original; // @[Interface.scala 259:14]
  wire [7:0] fifoTailReg_byte_original_1 = fifoTailReg[15:8]; // @[Interface.scala 258:39]
  wire [7:0] _fifoTailReg_T_13 = wrReqData__bits_strb[1] ? rPause_byte_wdata_1 : fifoTailReg_byte_original_1; // @[Interface.scala 259:14]
  wire [7:0] fifoTailReg_byte_original_2 = fifoTailReg[23:16]; // @[Interface.scala 258:39]
  wire [7:0] _fifoTailReg_T_14 = wrReqData__bits_strb[2] ? rPause_byte_wdata_2 : fifoTailReg_byte_original_2; // @[Interface.scala 259:14]
  wire [7:0] fifoTailReg_byte_original_3 = fifoTailReg[31:24]; // @[Interface.scala 258:39]
  wire [7:0] _fifoTailReg_T_15 = wrReqData__bits_strb[3] ? rPause_byte_wdata_3 : fifoTailReg_byte_original_3; // @[Interface.scala 259:14]
  wire [7:0] fifoTailReg_byte_original_4 = fifoTailReg[39:32]; // @[Interface.scala 258:39]
  wire [7:0] _fifoTailReg_T_16 = wrReqData__bits_strb[4] ? rPause_byte_wdata_4 : fifoTailReg_byte_original_4; // @[Interface.scala 259:14]
  wire [7:0] fifoTailReg_byte_original_5 = fifoTailReg[47:40]; // @[Interface.scala 258:39]
  wire [7:0] _fifoTailReg_T_17 = wrReqData__bits_strb[5] ? rPause_byte_wdata_5 : fifoTailReg_byte_original_5; // @[Interface.scala 259:14]
  wire [7:0] fifoTailReg_byte_original_6 = fifoTailReg[55:48]; // @[Interface.scala 258:39]
  wire [7:0] _fifoTailReg_T_18 = wrReqData__bits_strb[6] ? rPause_byte_wdata_6 : fifoTailReg_byte_original_6; // @[Interface.scala 259:14]
  wire [7:0] fifoTailReg_byte_original_7 = fifoTailReg[63:56]; // @[Interface.scala 258:39]
  wire [7:0] _fifoTailReg_T_19 = wrReqData__bits_strb[7] ? rPause_byte_wdata_7 : fifoTailReg_byte_original_7; // @[Interface.scala 259:14]
  wire [63:0] _fifoTailReg_T_20 = {_fifoTailReg_T_19,_fifoTailReg_T_18,_fifoTailReg_T_17,_fifoTailReg_T_16,
    _fifoTailReg_T_15,_fifoTailReg_T_14,_fifoTailReg_T_13,_fifoTailReg_T_12}; // @[Interface.scala 262:7]
  wire [7:0] fifoHeadReg_byte_original = fifoHeadReg[7:0]; // @[Interface.scala 258:39]
  wire [7:0] _fifoHeadReg_T_12 = wrReqData__bits_strb[0] ? rPause_byte_wdata : fifoHeadReg_byte_original; // @[Interface.scala 259:14]
  wire [7:0] fifoHeadReg_byte_original_1 = fifoHeadReg[15:8]; // @[Interface.scala 258:39]
  wire [7:0] _fifoHeadReg_T_13 = wrReqData__bits_strb[1] ? rPause_byte_wdata_1 : fifoHeadReg_byte_original_1; // @[Interface.scala 259:14]
  wire [7:0] fifoHeadReg_byte_original_2 = fifoHeadReg[23:16]; // @[Interface.scala 258:39]
  wire [7:0] _fifoHeadReg_T_14 = wrReqData__bits_strb[2] ? rPause_byte_wdata_2 : fifoHeadReg_byte_original_2; // @[Interface.scala 259:14]
  wire [7:0] fifoHeadReg_byte_original_3 = fifoHeadReg[31:24]; // @[Interface.scala 258:39]
  wire [7:0] _fifoHeadReg_T_15 = wrReqData__bits_strb[3] ? rPause_byte_wdata_3 : fifoHeadReg_byte_original_3; // @[Interface.scala 259:14]
  wire [7:0] fifoHeadReg_byte_original_4 = fifoHeadReg[39:32]; // @[Interface.scala 258:39]
  wire [7:0] _fifoHeadReg_T_16 = wrReqData__bits_strb[4] ? rPause_byte_wdata_4 : fifoHeadReg_byte_original_4; // @[Interface.scala 259:14]
  wire [7:0] fifoHeadReg_byte_original_5 = fifoHeadReg[47:40]; // @[Interface.scala 258:39]
  wire [7:0] _fifoHeadReg_T_17 = wrReqData__bits_strb[5] ? rPause_byte_wdata_5 : fifoHeadReg_byte_original_5; // @[Interface.scala 259:14]
  wire [7:0] fifoHeadReg_byte_original_6 = fifoHeadReg[55:48]; // @[Interface.scala 258:39]
  wire [7:0] _fifoHeadReg_T_18 = wrReqData__bits_strb[6] ? rPause_byte_wdata_6 : fifoHeadReg_byte_original_6; // @[Interface.scala 259:14]
  wire [7:0] fifoHeadReg_byte_original_7 = fifoHeadReg[63:56]; // @[Interface.scala 258:39]
  wire [7:0] _fifoHeadReg_T_19 = wrReqData__bits_strb[7] ? rPause_byte_wdata_7 : fifoHeadReg_byte_original_7; // @[Interface.scala 259:14]
  wire [63:0] _fifoHeadReg_T_20 = {_fifoHeadReg_T_19,_fifoHeadReg_T_18,_fifoHeadReg_T_17,_fifoHeadReg_T_16,
    _fifoHeadReg_T_15,_fifoHeadReg_T_14,_fifoHeadReg_T_13,_fifoHeadReg_T_12}; // @[Interface.scala 262:7]
  wire [7:0] procInterrupt_byte_original = procInterrupt[7:0]; // @[Interface.scala 258:39]
  wire [7:0] _procInterrupt_T_8 = wrReqData__bits_strb[0] ? rPause_byte_wdata : procInterrupt_byte_original; // @[Interface.scala 259:14]
  wire [7:0] procInterrupt_byte_original_1 = procInterrupt[15:8]; // @[Interface.scala 258:39]
  wire [7:0] _procInterrupt_T_9 = wrReqData__bits_strb[1] ? rPause_byte_wdata_1 : procInterrupt_byte_original_1; // @[Interface.scala 259:14]
  wire [7:0] procInterrupt_byte_original_2 = procInterrupt[23:16]; // @[Interface.scala 258:39]
  wire [7:0] _procInterrupt_T_10 = wrReqData__bits_strb[2] ? rPause_byte_wdata_2 : procInterrupt_byte_original_2; // @[Interface.scala 259:14]
  wire [7:0] procInterrupt_byte_original_3 = procInterrupt[31:24]; // @[Interface.scala 258:39]
  wire [7:0] _procInterrupt_T_11 = wrReqData__bits_strb[3] ? rPause_byte_wdata_3 : procInterrupt_byte_original_3; // @[Interface.scala 259:14]
  wire [7:0] procInterrupt_byte_original_4 = procInterrupt[39:32]; // @[Interface.scala 258:39]
  wire [7:0] _procInterrupt_T_12 = wrReqData__bits_strb[4] ? rPause_byte_wdata_4 : procInterrupt_byte_original_4; // @[Interface.scala 259:14]
  wire [7:0] procInterrupt_byte_original_5 = procInterrupt[47:40]; // @[Interface.scala 258:39]
  wire [7:0] _procInterrupt_T_13 = wrReqData__bits_strb[5] ? rPause_byte_wdata_5 : procInterrupt_byte_original_5; // @[Interface.scala 259:14]
  wire [7:0] procInterrupt_byte_original_6 = procInterrupt[55:48]; // @[Interface.scala 258:39]
  wire [7:0] _procInterrupt_T_14 = wrReqData__bits_strb[6] ? rPause_byte_wdata_6 : procInterrupt_byte_original_6; // @[Interface.scala 259:14]
  wire [7:0] procInterrupt_byte_original_7 = procInterrupt[63:56]; // @[Interface.scala 258:39]
  wire [7:0] _procInterrupt_T_15 = wrReqData__bits_strb[7] ? rPause_byte_wdata_7 : procInterrupt_byte_original_7; // @[Interface.scala 259:14]
  wire [63:0] _procInterrupt_T_16 = {_procInterrupt_T_15,_procInterrupt_T_14,_procInterrupt_T_13,_procInterrupt_T_12,
    _procInterrupt_T_11,_procInterrupt_T_10,_procInterrupt_T_9,_procInterrupt_T_8}; // @[Interface.scala 262:7]
  wire [63:0] _GEN_170 = reset ? 64'h0 : _GEN_74; // @[virtualStealServer.scala 82:{44,44}]
  Queue rdReq__deq ( // @[Decoupled.scala 377:21]
    .clock(rdReq__deq_clock),
    .reset(rdReq__deq_reset),
    .io_enq_ready(rdReq__deq_io_enq_ready),
    .io_enq_valid(rdReq__deq_io_enq_valid),
    .io_enq_bits_addr(rdReq__deq_io_enq_bits_addr),
    .io_deq_ready(rdReq__deq_io_deq_ready),
    .io_deq_valid(rdReq__deq_io_deq_valid),
    .io_deq_bits_addr(rdReq__deq_io_deq_bits_addr)
  );
  Queue wrReq__deq ( // @[Decoupled.scala 377:21]
    .clock(wrReq__deq_clock),
    .reset(wrReq__deq_reset),
    .io_enq_ready(wrReq__deq_io_enq_ready),
    .io_enq_valid(wrReq__deq_io_enq_valid),
    .io_enq_bits_addr(wrReq__deq_io_enq_bits_addr),
    .io_deq_ready(wrReq__deq_io_deq_ready),
    .io_deq_valid(wrReq__deq_io_deq_valid),
    .io_deq_bits_addr(wrReq__deq_io_deq_bits_addr)
  );
  Queue_2 wrReqData__deq ( // @[Decoupled.scala 377:21]
    .clock(wrReqData__deq_clock),
    .reset(wrReqData__deq_reset),
    .io_enq_ready(wrReqData__deq_io_enq_ready),
    .io_enq_valid(wrReqData__deq_io_enq_valid),
    .io_enq_bits_data(wrReqData__deq_io_enq_bits_data),
    .io_enq_bits_strb(wrReqData__deq_io_enq_bits_strb),
    .io_deq_ready(wrReqData__deq_io_deq_ready),
    .io_deq_valid(wrReqData__deq_io_deq_valid),
    .io_deq_bits_data(wrReqData__deq_io_deq_bits_data),
    .io_deq_bits_strb(wrReqData__deq_io_deq_bits_strb)
  );
  Queue_3 taskQueueBuffer ( // @[virtualStealServer.scala 81:43]
    .clock(taskQueueBuffer_clock),
    .reset(taskQueueBuffer_reset),
    .io_enq_ready(taskQueueBuffer_io_enq_ready),
    .io_enq_valid(taskQueueBuffer_io_enq_valid),
    .io_enq_bits(taskQueueBuffer_io_enq_bits),
    .io_deq_ready(taskQueueBuffer_io_deq_ready),
    .io_deq_valid(taskQueueBuffer_io_deq_valid),
    .io_deq_bits(taskQueueBuffer_io_deq_bits),
    .io_count(taskQueueBuffer_io_count)
  );
  assign io_connNetwork_ctrl_serveStealReq_valid = _T_29 ? 1'h0 : _GEN_122; // @[virtualStealServer.scala 309:40 293:45]
  assign io_connNetwork_data_availableTask_ready = stateReg == 4'h2; // @[virtualStealServer.scala 309:19]
  assign io_connNetwork_data_qOutTask_valid = _T_29 ? 1'h0 : _GEN_121; // @[virtualStealServer.scala 309:40 289:45]
  assign io_connNetwork_data_qOutTask_bits = taskQueueBuffer_io_deq_bits; // @[virtualStealServer.scala 275:45]
  assign io_axi_mgmt_ARREADY = rdReq__deq_io_enq_ready; // @[Decoupled.scala 381:17 RegisterBlock.scala 60:19]
  assign io_axi_mgmt_RVALID = rdReq__valid & io_axi_mgmt_RREADY; // @[RegisterBlock.scala 210:44]
  assign io_axi_mgmt_RDATA = 6'h28 == rdAddr ? procInterrupt : _GEN_147; // @[RegisterBlock.scala 224:38 225:16]
  assign io_axi_mgmt_AWREADY = wrReq__deq_io_enq_ready; // @[Decoupled.scala 381:17 RegisterBlock.scala 60:19]
  assign io_axi_mgmt_WREADY = wrReqData__deq_io_enq_ready; // @[Decoupled.scala 381:17 RegisterBlock.scala 60:19]
  assign io_axi_mgmt_BVALID = wrReq__valid & wrReqData__valid & io_axi_mgmt_BREADY; // @[RegisterBlock.scala 241:63]
  assign io_read_address_valid = _T_29 ? 1'h0 : _GEN_115; // @[virtualStealServer.scala 309:40 280:45]
  assign io_read_address_bits = _GEN_133[63:0];
  assign io_read_data_ready = _T_29 ? 1'h0 : _GEN_118; // @[virtualStealServer.scala 309:40 282:45]
  assign io_read_burst_len = _GEN_134[3:0];
  assign io_write_address_valid = _T_29 ? 1'h0 : _T_34; // @[virtualStealServer.scala 309:40 283:45]
  assign io_write_address_bits = _GEN_127[63:0];
  assign io_write_data_valid = _T_29 ? 1'h0 : _GEN_112; // @[virtualStealServer.scala 309:40 285:45]
  assign io_write_data_bits = taskQueueBuffer_io_deq_bits; // @[virtualStealServer.scala 276:45]
  assign io_write_burst_len = _T_29 ? 4'h0 : _GEN_111; // @[virtualStealServer.scala 309:40 302:45]
  assign io_write_last = _T_29 ? 1'h0 : _GEN_114; // @[virtualStealServer.scala 309:40 303:45]
  assign rdReq__deq_clock = clock;
  assign rdReq__deq_reset = reset;
  assign rdReq__deq_io_enq_valid = io_axi_mgmt_ARVALID; // @[RegisterBlock.scala 60:19 virtualStealServer.scala 62:20]
  assign rdReq__deq_io_enq_bits_addr = io_axi_mgmt_ARADDR; // @[RegisterBlock.scala 60:19 virtualStealServer.scala 62:20]
  assign rdReq__deq_io_deq_ready = rdReq__valid & io_axi_mgmt_RREADY; // @[RegisterBlock.scala 210:44]
  assign wrReq__deq_clock = clock;
  assign wrReq__deq_reset = reset;
  assign wrReq__deq_io_enq_valid = io_axi_mgmt_AWVALID; // @[RegisterBlock.scala 60:19 virtualStealServer.scala 62:20]
  assign wrReq__deq_io_enq_bits_addr = io_axi_mgmt_AWADDR; // @[RegisterBlock.scala 60:19 virtualStealServer.scala 62:20]
  assign wrReq__deq_io_deq_ready = wrReq__valid & wrReqData__valid & io_axi_mgmt_BREADY; // @[RegisterBlock.scala 241:63]
  assign wrReqData__deq_clock = clock;
  assign wrReqData__deq_reset = reset;
  assign wrReqData__deq_io_enq_valid = io_axi_mgmt_WVALID; // @[RegisterBlock.scala 60:19 virtualStealServer.scala 62:20]
  assign wrReqData__deq_io_enq_bits_data = io_axi_mgmt_WDATA; // @[RegisterBlock.scala 60:19 virtualStealServer.scala 62:20]
  assign wrReqData__deq_io_enq_bits_strb = io_axi_mgmt_WSTRB; // @[RegisterBlock.scala 60:19 virtualStealServer.scala 62:20]
  assign wrReqData__deq_io_deq_ready = wrReq__valid & wrReqData__valid & io_axi_mgmt_BREADY; // @[RegisterBlock.scala 241:63]
  assign taskQueueBuffer_clock = clock;
  assign taskQueueBuffer_reset = reset;
  assign taskQueueBuffer_io_enq_valid = _T_29 ? io_connNetwork_data_availableTask_valid : _GEN_120; // @[virtualStealServer.scala 309:40 313:49]
  assign taskQueueBuffer_io_enq_bits = _T_29 ? io_connNetwork_data_availableTask_bits : _GEN_119; // @[virtualStealServer.scala 309:40 311:49]
  assign taskQueueBuffer_io_deq_ready = _T_29 ? 1'h0 : _GEN_113; // @[virtualStealServer.scala 309:40 299:45]
  always @(posedge clock) begin
    if (reset) begin // @[virtualStealServer.scala 65:44]
      rAddr <= 64'h0; // @[virtualStealServer.scala 65:44]
    end else if (wrReq) begin // @[virtualStealServer.scala 388:27]
      if (6'h8 == wrAddr) begin // @[RegisterBlock.scala 252:38]
        rAddr <= _rAddr_T_16; // @[RegisterBlock.scala 118:11]
      end
    end
    if (reset) begin // @[virtualStealServer.scala 66:44]
      rPause <= 64'h0; // @[virtualStealServer.scala 66:44]
    end else if (wrReq) begin // @[virtualStealServer.scala 388:27]
      if (6'h0 == wrAddr) begin // @[RegisterBlock.scala 252:38]
        rPause <= _rPause_T_16; // @[RegisterBlock.scala 118:11]
      end else begin
        rPause <= _GEN_73;
      end
    end else begin
      rPause <= _GEN_73;
    end
    if (reset) begin // @[virtualStealServer.scala 67:44]
      procInterrupt <= 64'h0; // @[virtualStealServer.scala 67:44]
    end else if (wrReq) begin // @[virtualStealServer.scala 388:27]
      if (6'h28 == wrAddr) begin // @[RegisterBlock.scala 252:38]
        procInterrupt <= _procInterrupt_T_16; // @[RegisterBlock.scala 118:11]
      end
    end
    if (reset) begin // @[virtualStealServer.scala 68:44]
      maxLength <= 64'h0; // @[virtualStealServer.scala 68:44]
    end else if (wrReq) begin // @[virtualStealServer.scala 388:27]
      if (6'h10 == wrAddr) begin // @[RegisterBlock.scala 252:38]
        maxLength <= _maxLength_T_16; // @[RegisterBlock.scala 118:11]
      end
    end
    if (reset) begin // @[virtualStealServer.scala 69:44]
      stateReg <= 4'h0; // @[virtualStealServer.scala 69:44]
    end else if (stateReg == 4'h0) begin // @[virtualStealServer.scala 130:34]
      if (currLen == maxLength & networkCongested | maxLength < _T_15) begin // @[virtualStealServer.scala 132:90]
        stateReg <= 4'h9; // @[virtualStealServer.scala 134:22]
      end else if (networkCongested & taskQueueBuffer_io_count == 5'h10) begin // @[virtualStealServer.scala 137:74]
        stateReg <= 4'h4; // @[virtualStealServer.scala 139:22]
      end else begin
        stateReg <= _GEN_10;
      end
    end else if (stateReg == 4'h2) begin // @[virtualStealServer.scala 160:46]
      if (taskQueueBuffer_io_count == 5'hf & io_connNetwork_data_availableTask_valid) begin // @[virtualStealServer.scala 162:91]
        stateReg <= 4'h4; // @[virtualStealServer.scala 164:22]
      end else begin
        stateReg <= _GEN_17;
      end
    end else if (stateReg == 4'h4) begin // @[virtualStealServer.scala 176:54]
      stateReg <= _GEN_19;
    end else begin
      stateReg <= _GEN_57;
    end
    if (reset) begin // @[virtualStealServer.scala 71:44]
      contentionCounter <= 64'h0; // @[virtualStealServer.scala 71:44]
    end else if (io_ntwDataUnitOccupancy & contentionCounter != 64'h42) begin // @[virtualStealServer.scala 97:60]
      contentionCounter <= _contentionCounter_T_1; // @[virtualStealServer.scala 98:31]
    end else if (_T_2 & ~io_ntwDataUnitOccupancy) begin // @[virtualStealServer.scala 100:50]
      contentionCounter <= _contentionCounter_T_3; // @[virtualStealServer.scala 101:31]
    end
    if (reset) begin // @[virtualStealServer.scala 73:44]
      networkCongested <= 1'h0; // @[virtualStealServer.scala 73:44]
    end else begin
      networkCongested <= _GEN_3;
    end
    if (reset) begin // @[virtualStealServer.scala 77:44]
      fifoTailReg <= 64'h0; // @[virtualStealServer.scala 77:44]
    end else if (wrReq) begin // @[virtualStealServer.scala 388:27]
      if (6'h18 == wrAddr) begin // @[RegisterBlock.scala 252:38]
        fifoTailReg <= _fifoTailReg_T_20; // @[RegisterBlock.scala 118:11]
      end else begin
        fifoTailReg <= _GEN_76;
      end
    end else begin
      fifoTailReg <= _GEN_76;
    end
    if (reset) begin // @[virtualStealServer.scala 78:44]
      fifoHeadReg <= 64'h0; // @[virtualStealServer.scala 78:44]
    end else if (wrReq) begin // @[virtualStealServer.scala 388:27]
      if (6'h20 == wrAddr) begin // @[RegisterBlock.scala 252:38]
        fifoHeadReg <= _fifoHeadReg_T_20; // @[RegisterBlock.scala 118:11]
      end else begin
        fifoHeadReg <= _GEN_77;
      end
    end else begin
      fifoHeadReg <= _GEN_77;
    end
    popOrPush <= reset | _GEN_75; // @[virtualStealServer.scala 79:{44,44}]
    memDataCounter <= _GEN_170[4:0]; // @[virtualStealServer.scala 82:{44,44}]
    if (reset) begin // @[virtualStealServer.scala 355:32]
      lengthHistroy <= 64'h0; // @[virtualStealServer.scala 355:32]
    end else if (fifoTailReg > fifoHeadReg) begin // @[virtualStealServer.scala 357:36]
      lengthHistroy <= currLen; // @[virtualStealServer.scala 360:23]
    end else if (fifoTailReg < fifoHeadReg) begin // @[virtualStealServer.scala 362:42]
      lengthHistroy <= currLen; // @[virtualStealServer.scala 365:23]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rdReq & ~reset & ~rdReq) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegisterBlock.scala:182 assert(rdReq)\n"); // @[RegisterBlock.scala 182:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~rdReq & (rdReq & ~reset)) begin
          $fatal; // @[RegisterBlock.scala 182:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (wrReq & _T_77 & ~wrReq) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegisterBlock.scala:198 assert(wrReq)\n"); // @[RegisterBlock.scala 198:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~wrReq & (wrReq & _T_77)) begin
          $fatal; // @[RegisterBlock.scala 198:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  rAddr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  rPause = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  procInterrupt = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  maxLength = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  stateReg = _RAND_4[3:0];
  _RAND_5 = {2{`RANDOM}};
  contentionCounter = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  networkCongested = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  fifoTailReg = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  fifoHeadReg = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  popOrPush = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  memDataCounter = _RAND_10[4:0];
  _RAND_11 = {2{`RANDOM}};
  lengthHistroy = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module readyValidMem(
  input          clock,
  input          reset,
  output         io_read_address_ready,
  input          io_read_address_valid,
  input  [63:0]  io_read_address_bits,
  input          io_read_data_ready,
  output         io_read_data_valid,
  output [255:0] io_read_data_bits,
  output         io_write_address_ready,
  input          io_write_address_valid,
  input  [63:0]  io_write_address_bits,
  output         io_write_data_ready,
  input          io_write_data_valid,
  input  [255:0] io_write_data_bits,
  input  [3:0]   io_writeBurst_len,
  input          io_writeBurst_last,
  input  [3:0]   io_readBurst_len,
  input          axi_ARREADY,
  output         axi_ARVALID,
  output [63:0]  axi_ARADDR,
  output [7:0]   axi_ARLEN,
  output         axi_RREADY,
  input          axi_RVALID,
  input  [255:0] axi_RDATA,
  input          axi_AWREADY,
  output         axi_AWVALID,
  output [63:0]  axi_AWADDR,
  output [7:0]   axi_AWLEN,
  input          axi_WREADY,
  output         axi_WVALID,
  output [255:0] axi_WDATA,
  output         axi_WLAST,
  input          axi_BVALID
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  writeHandshakeDetector; // @[readyValidMem.scala 49:39]
  wire  _T_1 = ~writeHandshakeDetector; // @[readyValidMem.scala 81:58]
  wire  _GEN_0 = io_writeBurst_last | writeHandshakeDetector; // @[readyValidMem.scala 84:45 85:34 49:39]
  assign io_read_address_ready = axi_ARREADY; // @[readyValidMem.scala 155:31]
  assign io_read_data_valid = axi_RVALID; // @[readyValidMem.scala 171:31]
  assign io_read_data_bits = axi_RDATA; // @[readyValidMem.scala 172:31]
  assign io_write_address_ready = axi_AWREADY; // @[readyValidMem.scala 143:32]
  assign io_write_data_ready = axi_WREADY & _T_1; // @[readyValidMem.scala 94:53]
  assign axi_ARVALID = io_read_address_valid; // @[readyValidMem.scala 153:31]
  assign axi_ARADDR = io_read_address_bits; // @[readyValidMem.scala 154:31]
  assign axi_ARLEN = {{4'd0}, io_readBurst_len}; // @[readyValidMem.scala 158:33]
  assign axi_RREADY = io_read_data_ready; // @[readyValidMem.scala 169:31]
  assign axi_AWVALID = io_write_address_valid; // @[readyValidMem.scala 116:28]
  assign axi_AWADDR = io_write_address_bits; // @[readyValidMem.scala 117:28]
  assign axi_AWLEN = {{4'd0}, io_writeBurst_len}; // @[readyValidMem.scala 120:30]
  assign axi_WVALID = io_write_data_valid & axi_WREADY & ~writeHandshakeDetector; // @[readyValidMem.scala 81:55]
  assign axi_WDATA = io_write_data_bits; // @[readyValidMem.scala 130:28]
  assign axi_WLAST = io_writeBurst_last; // @[readyValidMem.scala 134:30]
  always @(posedge clock) begin
    if (reset) begin // @[readyValidMem.scala 49:39]
      writeHandshakeDetector <= 1'h0; // @[readyValidMem.scala 49:39]
    end else if (io_write_data_valid & axi_WREADY & ~writeHandshakeDetector) begin // @[readyValidMem.scala 81:82]
      writeHandshakeDetector <= _GEN_0;
    end else if (axi_BVALID) begin // @[readyValidMem.scala 88:34]
      writeHandshakeDetector <= 1'h0; // @[readyValidMem.scala 90:32]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeHandshakeDetector = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module stealSide(
  input          clock,
  input          reset,
  output         io_axi_mgmt_vss_0_ARREADY,
  input          io_axi_mgmt_vss_0_ARVALID,
  input  [5:0]   io_axi_mgmt_vss_0_ARADDR,
  input          io_axi_mgmt_vss_0_RREADY,
  output         io_axi_mgmt_vss_0_RVALID,
  output [63:0]  io_axi_mgmt_vss_0_RDATA,
  output         io_axi_mgmt_vss_0_AWREADY,
  input          io_axi_mgmt_vss_0_AWVALID,
  input  [5:0]   io_axi_mgmt_vss_0_AWADDR,
  output         io_axi_mgmt_vss_0_WREADY,
  input          io_axi_mgmt_vss_0_WVALID,
  input  [63:0]  io_axi_mgmt_vss_0_WDATA,
  input  [7:0]   io_axi_mgmt_vss_0_WSTRB,
  input          io_axi_mgmt_vss_0_BREADY,
  output         io_axi_mgmt_vss_0_BVALID,
  input          io_vss_axi_full_0_ARREADY,
  output         io_vss_axi_full_0_ARVALID,
  output [63:0]  io_vss_axi_full_0_ARADDR,
  output [7:0]   io_vss_axi_full_0_ARLEN,
  output         io_vss_axi_full_0_RREADY,
  input          io_vss_axi_full_0_RVALID,
  input  [255:0] io_vss_axi_full_0_RDATA,
  input          io_vss_axi_full_0_AWREADY,
  output         io_vss_axi_full_0_AWVALID,
  output [63:0]  io_vss_axi_full_0_AWADDR,
  output [7:0]   io_vss_axi_full_0_AWLEN,
  input          io_vss_axi_full_0_WREADY,
  output         io_vss_axi_full_0_WVALID,
  output [255:0] io_vss_axi_full_0_WDATA,
  output         io_vss_axi_full_0_WLAST,
  input          io_vss_axi_full_0_BVALID,
  input          io_taskOut_0_TREADY,
  output         io_taskOut_0_TVALID,
  output [255:0] io_taskOut_0_TDATA,
  input          io_taskOut_1_TREADY,
  output         io_taskOut_1_TVALID,
  output [255:0] io_taskOut_1_TDATA,
  input          io_taskOut_2_TREADY,
  output         io_taskOut_2_TVALID,
  output [255:0] io_taskOut_2_TDATA,
  input          io_taskOut_3_TREADY,
  output         io_taskOut_3_TVALID,
  output [255:0] io_taskOut_3_TDATA,
  input          io_taskOut_4_TREADY,
  output         io_taskOut_4_TVALID,
  output [255:0] io_taskOut_4_TDATA,
  input          io_taskOut_5_TREADY,
  output         io_taskOut_5_TVALID,
  output [255:0] io_taskOut_5_TDATA,
  input          io_taskOut_6_TREADY,
  output         io_taskOut_6_TVALID,
  output [255:0] io_taskOut_6_TDATA,
  input          io_taskOut_7_TREADY,
  output         io_taskOut_7_TVALID,
  output [255:0] io_taskOut_7_TDATA,
  input          io_taskOut_8_TREADY,
  output         io_taskOut_8_TVALID,
  output [255:0] io_taskOut_8_TDATA,
  input          io_taskOut_9_TREADY,
  output         io_taskOut_9_TVALID,
  output [255:0] io_taskOut_9_TDATA,
  input          io_taskOut_10_TREADY,
  output         io_taskOut_10_TVALID,
  output [255:0] io_taskOut_10_TDATA,
  input          io_taskOut_11_TREADY,
  output         io_taskOut_11_TVALID,
  output [255:0] io_taskOut_11_TDATA,
  input          io_taskOut_12_TREADY,
  output         io_taskOut_12_TVALID,
  output [255:0] io_taskOut_12_TDATA,
  input          io_taskOut_13_TREADY,
  output         io_taskOut_13_TVALID,
  output [255:0] io_taskOut_13_TDATA,
  input          io_taskOut_14_TREADY,
  output         io_taskOut_14_TVALID,
  output [255:0] io_taskOut_14_TDATA,
  input          io_taskOut_15_TREADY,
  output         io_taskOut_15_TVALID,
  output [255:0] io_taskOut_15_TDATA,
  input          io_taskOut_16_TREADY,
  output         io_taskOut_16_TVALID,
  output [255:0] io_taskOut_16_TDATA,
  input          io_taskOut_17_TREADY,
  output         io_taskOut_17_TVALID,
  output [255:0] io_taskOut_17_TDATA,
  input          io_taskOut_18_TREADY,
  output         io_taskOut_18_TVALID,
  output [255:0] io_taskOut_18_TDATA,
  input          io_taskOut_19_TREADY,
  output         io_taskOut_19_TVALID,
  output [255:0] io_taskOut_19_TDATA,
  input          io_taskOut_20_TREADY,
  output         io_taskOut_20_TVALID,
  output [255:0] io_taskOut_20_TDATA,
  input          io_taskOut_21_TREADY,
  output         io_taskOut_21_TVALID,
  output [255:0] io_taskOut_21_TDATA,
  input          io_taskOut_22_TREADY,
  output         io_taskOut_22_TVALID,
  output [255:0] io_taskOut_22_TDATA,
  input          io_taskOut_23_TREADY,
  output         io_taskOut_23_TVALID,
  output [255:0] io_taskOut_23_TDATA,
  input          io_taskOut_24_TREADY,
  output         io_taskOut_24_TVALID,
  output [255:0] io_taskOut_24_TDATA,
  input          io_taskOut_25_TREADY,
  output         io_taskOut_25_TVALID,
  output [255:0] io_taskOut_25_TDATA,
  input          io_taskOut_26_TREADY,
  output         io_taskOut_26_TVALID,
  output [255:0] io_taskOut_26_TDATA,
  input          io_taskOut_27_TREADY,
  output         io_taskOut_27_TVALID,
  output [255:0] io_taskOut_27_TDATA,
  input          io_taskOut_28_TREADY,
  output         io_taskOut_28_TVALID,
  output [255:0] io_taskOut_28_TDATA,
  input          io_taskOut_29_TREADY,
  output         io_taskOut_29_TVALID,
  output [255:0] io_taskOut_29_TDATA,
  input          io_taskOut_30_TREADY,
  output         io_taskOut_30_TVALID,
  output [255:0] io_taskOut_30_TDATA,
  input          io_taskOut_31_TREADY,
  output         io_taskOut_31_TVALID,
  output [255:0] io_taskOut_31_TDATA,
  input          io_taskOut_32_TREADY,
  output         io_taskOut_32_TVALID,
  output [255:0] io_taskOut_32_TDATA,
  input          io_taskOut_33_TREADY,
  output         io_taskOut_33_TVALID,
  output [255:0] io_taskOut_33_TDATA,
  input          io_taskOut_34_TREADY,
  output         io_taskOut_34_TVALID,
  output [255:0] io_taskOut_34_TDATA,
  input          io_taskOut_35_TREADY,
  output         io_taskOut_35_TVALID,
  output [255:0] io_taskOut_35_TDATA,
  input          io_taskOut_36_TREADY,
  output         io_taskOut_36_TVALID,
  output [255:0] io_taskOut_36_TDATA,
  input          io_taskOut_37_TREADY,
  output         io_taskOut_37_TVALID,
  output [255:0] io_taskOut_37_TDATA,
  input          io_taskOut_38_TREADY,
  output         io_taskOut_38_TVALID,
  output [255:0] io_taskOut_38_TDATA,
  input          io_taskOut_39_TREADY,
  output         io_taskOut_39_TVALID,
  output [255:0] io_taskOut_39_TDATA,
  input          io_taskOut_40_TREADY,
  output         io_taskOut_40_TVALID,
  output [255:0] io_taskOut_40_TDATA,
  input          io_taskOut_41_TREADY,
  output         io_taskOut_41_TVALID,
  output [255:0] io_taskOut_41_TDATA,
  input          io_taskOut_42_TREADY,
  output         io_taskOut_42_TVALID,
  output [255:0] io_taskOut_42_TDATA,
  input          io_taskOut_43_TREADY,
  output         io_taskOut_43_TVALID,
  output [255:0] io_taskOut_43_TDATA,
  input          io_taskOut_44_TREADY,
  output         io_taskOut_44_TVALID,
  output [255:0] io_taskOut_44_TDATA,
  input          io_taskOut_45_TREADY,
  output         io_taskOut_45_TVALID,
  output [255:0] io_taskOut_45_TDATA,
  input          io_taskOut_46_TREADY,
  output         io_taskOut_46_TVALID,
  output [255:0] io_taskOut_46_TDATA,
  input          io_taskOut_47_TREADY,
  output         io_taskOut_47_TVALID,
  output [255:0] io_taskOut_47_TDATA,
  input          io_taskOut_48_TREADY,
  output         io_taskOut_48_TVALID,
  output [255:0] io_taskOut_48_TDATA,
  input          io_taskOut_49_TREADY,
  output         io_taskOut_49_TVALID,
  output [255:0] io_taskOut_49_TDATA,
  input          io_taskOut_50_TREADY,
  output         io_taskOut_50_TVALID,
  output [255:0] io_taskOut_50_TDATA,
  input          io_taskOut_51_TREADY,
  output         io_taskOut_51_TVALID,
  output [255:0] io_taskOut_51_TDATA,
  input          io_taskOut_52_TREADY,
  output         io_taskOut_52_TVALID,
  output [255:0] io_taskOut_52_TDATA,
  input          io_taskOut_53_TREADY,
  output         io_taskOut_53_TVALID,
  output [255:0] io_taskOut_53_TDATA,
  input          io_taskOut_54_TREADY,
  output         io_taskOut_54_TVALID,
  output [255:0] io_taskOut_54_TDATA,
  input          io_taskOut_55_TREADY,
  output         io_taskOut_55_TVALID,
  output [255:0] io_taskOut_55_TDATA,
  input          io_taskOut_56_TREADY,
  output         io_taskOut_56_TVALID,
  output [255:0] io_taskOut_56_TDATA,
  input          io_taskOut_57_TREADY,
  output         io_taskOut_57_TVALID,
  output [255:0] io_taskOut_57_TDATA,
  input          io_taskOut_58_TREADY,
  output         io_taskOut_58_TVALID,
  output [255:0] io_taskOut_58_TDATA,
  input          io_taskOut_59_TREADY,
  output         io_taskOut_59_TVALID,
  output [255:0] io_taskOut_59_TDATA,
  input          io_taskOut_60_TREADY,
  output         io_taskOut_60_TVALID,
  output [255:0] io_taskOut_60_TDATA,
  input          io_taskOut_61_TREADY,
  output         io_taskOut_61_TVALID,
  output [255:0] io_taskOut_61_TDATA,
  input          io_taskOut_62_TREADY,
  output         io_taskOut_62_TVALID,
  output [255:0] io_taskOut_62_TDATA,
  input          io_taskOut_63_TREADY,
  output         io_taskOut_63_TVALID,
  output [255:0] io_taskOut_63_TDATA,
  output         io_taskIn_0_TREADY,
  input          io_taskIn_0_TVALID,
  input  [255:0] io_taskIn_0_TDATA,
  output         io_taskIn_1_TREADY,
  input          io_taskIn_1_TVALID,
  input  [255:0] io_taskIn_1_TDATA,
  output         io_taskIn_2_TREADY,
  input          io_taskIn_2_TVALID,
  input  [255:0] io_taskIn_2_TDATA,
  output         io_taskIn_3_TREADY,
  input          io_taskIn_3_TVALID,
  input  [255:0] io_taskIn_3_TDATA,
  output         io_taskIn_4_TREADY,
  input          io_taskIn_4_TVALID,
  input  [255:0] io_taskIn_4_TDATA,
  output         io_taskIn_5_TREADY,
  input          io_taskIn_5_TVALID,
  input  [255:0] io_taskIn_5_TDATA,
  output         io_taskIn_6_TREADY,
  input          io_taskIn_6_TVALID,
  input  [255:0] io_taskIn_6_TDATA,
  output         io_taskIn_7_TREADY,
  input          io_taskIn_7_TVALID,
  input  [255:0] io_taskIn_7_TDATA,
  output         io_taskIn_8_TREADY,
  input          io_taskIn_8_TVALID,
  input  [255:0] io_taskIn_8_TDATA,
  output         io_taskIn_9_TREADY,
  input          io_taskIn_9_TVALID,
  input  [255:0] io_taskIn_9_TDATA,
  output         io_taskIn_10_TREADY,
  input          io_taskIn_10_TVALID,
  input  [255:0] io_taskIn_10_TDATA,
  output         io_taskIn_11_TREADY,
  input          io_taskIn_11_TVALID,
  input  [255:0] io_taskIn_11_TDATA,
  output         io_taskIn_12_TREADY,
  input          io_taskIn_12_TVALID,
  input  [255:0] io_taskIn_12_TDATA,
  output         io_taskIn_13_TREADY,
  input          io_taskIn_13_TVALID,
  input  [255:0] io_taskIn_13_TDATA,
  output         io_taskIn_14_TREADY,
  input          io_taskIn_14_TVALID,
  input  [255:0] io_taskIn_14_TDATA,
  output         io_taskIn_15_TREADY,
  input          io_taskIn_15_TVALID,
  input  [255:0] io_taskIn_15_TDATA,
  output         io_taskIn_16_TREADY,
  input          io_taskIn_16_TVALID,
  input  [255:0] io_taskIn_16_TDATA,
  output         io_taskIn_17_TREADY,
  input          io_taskIn_17_TVALID,
  input  [255:0] io_taskIn_17_TDATA,
  output         io_taskIn_18_TREADY,
  input          io_taskIn_18_TVALID,
  input  [255:0] io_taskIn_18_TDATA,
  output         io_taskIn_19_TREADY,
  input          io_taskIn_19_TVALID,
  input  [255:0] io_taskIn_19_TDATA,
  output         io_taskIn_20_TREADY,
  input          io_taskIn_20_TVALID,
  input  [255:0] io_taskIn_20_TDATA,
  output         io_taskIn_21_TREADY,
  input          io_taskIn_21_TVALID,
  input  [255:0] io_taskIn_21_TDATA,
  output         io_taskIn_22_TREADY,
  input          io_taskIn_22_TVALID,
  input  [255:0] io_taskIn_22_TDATA,
  output         io_taskIn_23_TREADY,
  input          io_taskIn_23_TVALID,
  input  [255:0] io_taskIn_23_TDATA,
  output         io_taskIn_24_TREADY,
  input          io_taskIn_24_TVALID,
  input  [255:0] io_taskIn_24_TDATA,
  output         io_taskIn_25_TREADY,
  input          io_taskIn_25_TVALID,
  input  [255:0] io_taskIn_25_TDATA,
  output         io_taskIn_26_TREADY,
  input          io_taskIn_26_TVALID,
  input  [255:0] io_taskIn_26_TDATA,
  output         io_taskIn_27_TREADY,
  input          io_taskIn_27_TVALID,
  input  [255:0] io_taskIn_27_TDATA,
  output         io_taskIn_28_TREADY,
  input          io_taskIn_28_TVALID,
  input  [255:0] io_taskIn_28_TDATA,
  output         io_taskIn_29_TREADY,
  input          io_taskIn_29_TVALID,
  input  [255:0] io_taskIn_29_TDATA,
  output         io_taskIn_30_TREADY,
  input          io_taskIn_30_TVALID,
  input  [255:0] io_taskIn_30_TDATA,
  output         io_taskIn_31_TREADY,
  input          io_taskIn_31_TVALID,
  input  [255:0] io_taskIn_31_TDATA,
  output         io_taskIn_32_TREADY,
  input          io_taskIn_32_TVALID,
  input  [255:0] io_taskIn_32_TDATA,
  output         io_taskIn_33_TREADY,
  input          io_taskIn_33_TVALID,
  input  [255:0] io_taskIn_33_TDATA,
  output         io_taskIn_34_TREADY,
  input          io_taskIn_34_TVALID,
  input  [255:0] io_taskIn_34_TDATA,
  output         io_taskIn_35_TREADY,
  input          io_taskIn_35_TVALID,
  input  [255:0] io_taskIn_35_TDATA,
  output         io_taskIn_36_TREADY,
  input          io_taskIn_36_TVALID,
  input  [255:0] io_taskIn_36_TDATA,
  output         io_taskIn_37_TREADY,
  input          io_taskIn_37_TVALID,
  input  [255:0] io_taskIn_37_TDATA,
  output         io_taskIn_38_TREADY,
  input          io_taskIn_38_TVALID,
  input  [255:0] io_taskIn_38_TDATA,
  output         io_taskIn_39_TREADY,
  input          io_taskIn_39_TVALID,
  input  [255:0] io_taskIn_39_TDATA,
  output         io_taskIn_40_TREADY,
  input          io_taskIn_40_TVALID,
  input  [255:0] io_taskIn_40_TDATA,
  output         io_taskIn_41_TREADY,
  input          io_taskIn_41_TVALID,
  input  [255:0] io_taskIn_41_TDATA,
  output         io_taskIn_42_TREADY,
  input          io_taskIn_42_TVALID,
  input  [255:0] io_taskIn_42_TDATA,
  output         io_taskIn_43_TREADY,
  input          io_taskIn_43_TVALID,
  input  [255:0] io_taskIn_43_TDATA,
  output         io_taskIn_44_TREADY,
  input          io_taskIn_44_TVALID,
  input  [255:0] io_taskIn_44_TDATA,
  output         io_taskIn_45_TREADY,
  input          io_taskIn_45_TVALID,
  input  [255:0] io_taskIn_45_TDATA,
  output         io_taskIn_46_TREADY,
  input          io_taskIn_46_TVALID,
  input  [255:0] io_taskIn_46_TDATA,
  output         io_taskIn_47_TREADY,
  input          io_taskIn_47_TVALID,
  input  [255:0] io_taskIn_47_TDATA,
  output         io_taskIn_48_TREADY,
  input          io_taskIn_48_TVALID,
  input  [255:0] io_taskIn_48_TDATA,
  output         io_taskIn_49_TREADY,
  input          io_taskIn_49_TVALID,
  input  [255:0] io_taskIn_49_TDATA,
  output         io_taskIn_50_TREADY,
  input          io_taskIn_50_TVALID,
  input  [255:0] io_taskIn_50_TDATA,
  output         io_taskIn_51_TREADY,
  input          io_taskIn_51_TVALID,
  input  [255:0] io_taskIn_51_TDATA,
  output         io_taskIn_52_TREADY,
  input          io_taskIn_52_TVALID,
  input  [255:0] io_taskIn_52_TDATA,
  output         io_taskIn_53_TREADY,
  input          io_taskIn_53_TVALID,
  input  [255:0] io_taskIn_53_TDATA,
  output         io_taskIn_54_TREADY,
  input          io_taskIn_54_TVALID,
  input  [255:0] io_taskIn_54_TDATA,
  output         io_taskIn_55_TREADY,
  input          io_taskIn_55_TVALID,
  input  [255:0] io_taskIn_55_TDATA,
  output         io_taskIn_56_TREADY,
  input          io_taskIn_56_TVALID,
  input  [255:0] io_taskIn_56_TDATA,
  output         io_taskIn_57_TREADY,
  input          io_taskIn_57_TVALID,
  input  [255:0] io_taskIn_57_TDATA,
  output         io_taskIn_58_TREADY,
  input          io_taskIn_58_TVALID,
  input  [255:0] io_taskIn_58_TDATA,
  output         io_taskIn_59_TREADY,
  input          io_taskIn_59_TVALID,
  input  [255:0] io_taskIn_59_TDATA,
  output         io_taskIn_60_TREADY,
  input          io_taskIn_60_TVALID,
  input  [255:0] io_taskIn_60_TDATA,
  output         io_taskIn_61_TREADY,
  input          io_taskIn_61_TVALID,
  input  [255:0] io_taskIn_61_TDATA,
  output         io_taskIn_62_TREADY,
  input          io_taskIn_62_TVALID,
  input  [255:0] io_taskIn_62_TDATA,
  output         io_taskIn_63_TREADY,
  input          io_taskIn_63_TVALID,
  input  [255:0] io_taskIn_63_TDATA,
  output         connSyncSide_0_ctrl_serveStealReq_ready,
  input          connSyncSide_0_ctrl_serveStealReq_valid,
  output         connSyncSide_0_data_qOutTask_ready,
  input          connSyncSide_0_data_qOutTask_valid,
  input  [255:0] connSyncSide_0_data_qOutTask_bits,
  output         connSyncSide_1_ctrl_serveStealReq_ready,
  input          connSyncSide_1_ctrl_serveStealReq_valid,
  output         connSyncSide_1_data_qOutTask_ready,
  input          connSyncSide_1_data_qOutTask_valid,
  input  [255:0] connSyncSide_1_data_qOutTask_bits
);
  wire  stealNW_TQ_clock; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_reset; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_0_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_0_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_0_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_0_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_0_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_0_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_1_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_1_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_1_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_1_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_1_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_1_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_2_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_2_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_2_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_2_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_2_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_2_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_3_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_3_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_3_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_3_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_3_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_3_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_4_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_4_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_4_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_4_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_4_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_4_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_5_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_5_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_5_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_5_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_5_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_5_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_6_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_6_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_6_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_6_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_6_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_6_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_7_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_7_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_7_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_7_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_7_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_7_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_8_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_8_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_8_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_8_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_8_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_8_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_9_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_9_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_9_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_9_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_9_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_9_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_10_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_10_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_10_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_10_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_10_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_10_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_11_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_11_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_11_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_11_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_11_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_11_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_12_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_12_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_12_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_12_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_12_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_12_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_13_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_13_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_13_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_13_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_13_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_13_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_14_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_14_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_14_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_14_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_14_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_14_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_15_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_15_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_15_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_15_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_15_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_15_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_16_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_16_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_16_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_16_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_16_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_16_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_17_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_17_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_17_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_17_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_17_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_17_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_18_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_18_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_18_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_18_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_18_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_18_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_19_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_19_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_19_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_19_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_19_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_19_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_20_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_20_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_20_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_20_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_20_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_20_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_21_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_21_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_21_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_21_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_21_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_21_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_22_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_22_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_22_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_22_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_22_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_22_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_23_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_23_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_23_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_23_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_23_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_23_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_24_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_24_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_24_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_24_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_24_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_24_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_25_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_25_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_25_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_25_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_25_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_25_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_26_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_26_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_26_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_26_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_26_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_26_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_27_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_27_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_27_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_27_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_27_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_27_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_28_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_28_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_28_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_28_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_28_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_28_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_29_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_29_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_29_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_29_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_29_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_29_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_30_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_30_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_30_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_30_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_30_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_30_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_31_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_31_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_31_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_31_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_31_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_31_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_32_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_32_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_32_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_32_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_32_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_32_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_33_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_33_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_33_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_33_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_33_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_33_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_34_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_34_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_34_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_34_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_34_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_34_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_35_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_35_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_35_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_35_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_35_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_35_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_36_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_36_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_36_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_36_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_36_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_36_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_37_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_37_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_37_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_37_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_37_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_37_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_38_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_38_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_38_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_38_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_38_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_38_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_39_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_39_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_39_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_39_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_39_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_39_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_40_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_40_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_40_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_40_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_40_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_40_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_41_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_41_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_41_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_41_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_41_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_41_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_42_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_42_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_42_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_42_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_42_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_42_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_43_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_43_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_43_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_43_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_43_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_43_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_44_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_44_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_44_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_44_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_44_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_44_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_45_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_45_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_45_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_45_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_45_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_45_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_46_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_46_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_46_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_46_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_46_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_46_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_47_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_47_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_47_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_47_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_47_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_47_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_48_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_48_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_48_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_48_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_48_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_48_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_49_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_49_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_49_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_49_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_49_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_49_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_50_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_50_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_50_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_50_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_50_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_50_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_51_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_51_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_51_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_51_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_51_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_51_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_52_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_52_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_52_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_52_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_52_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_52_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_53_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_53_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_53_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_53_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_53_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_53_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_54_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_54_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_54_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_54_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_54_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_54_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_55_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_55_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_55_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_55_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_55_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_55_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_56_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_56_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_56_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_56_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_56_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_56_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_57_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_57_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_57_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_57_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_57_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_57_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_58_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_58_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_58_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_58_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_58_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_58_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_59_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_59_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_59_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_59_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_59_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_59_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_60_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_60_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_60_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_60_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_60_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_60_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_61_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_61_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_61_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_61_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_61_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_61_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_62_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_62_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_62_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_62_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_62_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_62_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_63_push_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_63_push_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_63_push_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_63_pop_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connPE_63_pop_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connPE_63_pop_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connVSS_0_ctrl_serveStealReq_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connVSS_0_ctrl_serveStealReq_valid; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connVSS_0_data_availableTask_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connVSS_0_data_availableTask_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connVSS_0_data_availableTask_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connVSS_0_data_qOutTask_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connVSS_0_data_qOutTask_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connVSS_0_data_qOutTask_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connVAS_0_ctrl_serveStealReq_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connVAS_0_ctrl_serveStealReq_valid; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connVAS_0_data_qOutTask_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connVAS_0_data_qOutTask_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connVAS_0_data_qOutTask_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connVAS_1_ctrl_serveStealReq_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connVAS_1_ctrl_serveStealReq_valid; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connVAS_1_data_qOutTask_ready; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_connVAS_1_data_qOutTask_valid; // @[stealSide.scala 55:28]
  wire [255:0] stealNW_TQ_io_connVAS_1_data_qOutTask_bits; // @[stealSide.scala 55:28]
  wire  stealNW_TQ_io_ntwDataUnitOccupancyVSS_0; // @[stealSide.scala 55:28]
  wire  virtualStealServers_0_clock; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_reset; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_connNetwork_ctrl_serveStealReq_ready; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_connNetwork_ctrl_serveStealReq_valid; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_connNetwork_data_availableTask_ready; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_connNetwork_data_availableTask_valid; // @[stealSide.scala 66:75]
  wire [255:0] virtualStealServers_0_io_connNetwork_data_availableTask_bits; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_connNetwork_data_qOutTask_ready; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_connNetwork_data_qOutTask_valid; // @[stealSide.scala 66:75]
  wire [255:0] virtualStealServers_0_io_connNetwork_data_qOutTask_bits; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_axi_mgmt_ARREADY; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_axi_mgmt_ARVALID; // @[stealSide.scala 66:75]
  wire [5:0] virtualStealServers_0_io_axi_mgmt_ARADDR; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_axi_mgmt_RREADY; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_axi_mgmt_RVALID; // @[stealSide.scala 66:75]
  wire [63:0] virtualStealServers_0_io_axi_mgmt_RDATA; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_axi_mgmt_AWREADY; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_axi_mgmt_AWVALID; // @[stealSide.scala 66:75]
  wire [5:0] virtualStealServers_0_io_axi_mgmt_AWADDR; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_axi_mgmt_WREADY; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_axi_mgmt_WVALID; // @[stealSide.scala 66:75]
  wire [63:0] virtualStealServers_0_io_axi_mgmt_WDATA; // @[stealSide.scala 66:75]
  wire [7:0] virtualStealServers_0_io_axi_mgmt_WSTRB; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_axi_mgmt_BREADY; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_axi_mgmt_BVALID; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_read_address_ready; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_read_address_valid; // @[stealSide.scala 66:75]
  wire [63:0] virtualStealServers_0_io_read_address_bits; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_read_data_ready; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_read_data_valid; // @[stealSide.scala 66:75]
  wire [255:0] virtualStealServers_0_io_read_data_bits; // @[stealSide.scala 66:75]
  wire [3:0] virtualStealServers_0_io_read_burst_len; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_write_address_ready; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_write_address_valid; // @[stealSide.scala 66:75]
  wire [63:0] virtualStealServers_0_io_write_address_bits; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_write_data_ready; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_write_data_valid; // @[stealSide.scala 66:75]
  wire [255:0] virtualStealServers_0_io_write_data_bits; // @[stealSide.scala 66:75]
  wire [3:0] virtualStealServers_0_io_write_burst_len; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_write_last; // @[stealSide.scala 66:75]
  wire  virtualStealServers_0_io_ntwDataUnitOccupancy; // @[stealSide.scala 66:75]
  wire  vssRvm_0_clock; // @[stealSide.scala 91:68]
  wire  vssRvm_0_reset; // @[stealSide.scala 91:68]
  wire  vssRvm_0_io_read_address_ready; // @[stealSide.scala 91:68]
  wire  vssRvm_0_io_read_address_valid; // @[stealSide.scala 91:68]
  wire [63:0] vssRvm_0_io_read_address_bits; // @[stealSide.scala 91:68]
  wire  vssRvm_0_io_read_data_ready; // @[stealSide.scala 91:68]
  wire  vssRvm_0_io_read_data_valid; // @[stealSide.scala 91:68]
  wire [255:0] vssRvm_0_io_read_data_bits; // @[stealSide.scala 91:68]
  wire  vssRvm_0_io_write_address_ready; // @[stealSide.scala 91:68]
  wire  vssRvm_0_io_write_address_valid; // @[stealSide.scala 91:68]
  wire [63:0] vssRvm_0_io_write_address_bits; // @[stealSide.scala 91:68]
  wire  vssRvm_0_io_write_data_ready; // @[stealSide.scala 91:68]
  wire  vssRvm_0_io_write_data_valid; // @[stealSide.scala 91:68]
  wire [255:0] vssRvm_0_io_write_data_bits; // @[stealSide.scala 91:68]
  wire [3:0] vssRvm_0_io_writeBurst_len; // @[stealSide.scala 91:68]
  wire  vssRvm_0_io_writeBurst_last; // @[stealSide.scala 91:68]
  wire [3:0] vssRvm_0_io_readBurst_len; // @[stealSide.scala 91:68]
  wire  vssRvm_0_axi_ARREADY; // @[stealSide.scala 91:68]
  wire  vssRvm_0_axi_ARVALID; // @[stealSide.scala 91:68]
  wire [63:0] vssRvm_0_axi_ARADDR; // @[stealSide.scala 91:68]
  wire [7:0] vssRvm_0_axi_ARLEN; // @[stealSide.scala 91:68]
  wire  vssRvm_0_axi_RREADY; // @[stealSide.scala 91:68]
  wire  vssRvm_0_axi_RVALID; // @[stealSide.scala 91:68]
  wire [255:0] vssRvm_0_axi_RDATA; // @[stealSide.scala 91:68]
  wire  vssRvm_0_axi_AWREADY; // @[stealSide.scala 91:68]
  wire  vssRvm_0_axi_AWVALID; // @[stealSide.scala 91:68]
  wire [63:0] vssRvm_0_axi_AWADDR; // @[stealSide.scala 91:68]
  wire [7:0] vssRvm_0_axi_AWLEN; // @[stealSide.scala 91:68]
  wire  vssRvm_0_axi_WREADY; // @[stealSide.scala 91:68]
  wire  vssRvm_0_axi_WVALID; // @[stealSide.scala 91:68]
  wire [255:0] vssRvm_0_axi_WDATA; // @[stealSide.scala 91:68]
  wire  vssRvm_0_axi_WLAST; // @[stealSide.scala 91:68]
  wire  vssRvm_0_axi_BVALID; // @[stealSide.scala 91:68]
  stealNW_TQ stealNW_TQ ( // @[stealSide.scala 55:28]
    .clock(stealNW_TQ_clock),
    .reset(stealNW_TQ_reset),
    .io_connPE_0_push_ready(stealNW_TQ_io_connPE_0_push_ready),
    .io_connPE_0_push_valid(stealNW_TQ_io_connPE_0_push_valid),
    .io_connPE_0_push_bits(stealNW_TQ_io_connPE_0_push_bits),
    .io_connPE_0_pop_ready(stealNW_TQ_io_connPE_0_pop_ready),
    .io_connPE_0_pop_valid(stealNW_TQ_io_connPE_0_pop_valid),
    .io_connPE_0_pop_bits(stealNW_TQ_io_connPE_0_pop_bits),
    .io_connPE_1_push_ready(stealNW_TQ_io_connPE_1_push_ready),
    .io_connPE_1_push_valid(stealNW_TQ_io_connPE_1_push_valid),
    .io_connPE_1_push_bits(stealNW_TQ_io_connPE_1_push_bits),
    .io_connPE_1_pop_ready(stealNW_TQ_io_connPE_1_pop_ready),
    .io_connPE_1_pop_valid(stealNW_TQ_io_connPE_1_pop_valid),
    .io_connPE_1_pop_bits(stealNW_TQ_io_connPE_1_pop_bits),
    .io_connPE_2_push_ready(stealNW_TQ_io_connPE_2_push_ready),
    .io_connPE_2_push_valid(stealNW_TQ_io_connPE_2_push_valid),
    .io_connPE_2_push_bits(stealNW_TQ_io_connPE_2_push_bits),
    .io_connPE_2_pop_ready(stealNW_TQ_io_connPE_2_pop_ready),
    .io_connPE_2_pop_valid(stealNW_TQ_io_connPE_2_pop_valid),
    .io_connPE_2_pop_bits(stealNW_TQ_io_connPE_2_pop_bits),
    .io_connPE_3_push_ready(stealNW_TQ_io_connPE_3_push_ready),
    .io_connPE_3_push_valid(stealNW_TQ_io_connPE_3_push_valid),
    .io_connPE_3_push_bits(stealNW_TQ_io_connPE_3_push_bits),
    .io_connPE_3_pop_ready(stealNW_TQ_io_connPE_3_pop_ready),
    .io_connPE_3_pop_valid(stealNW_TQ_io_connPE_3_pop_valid),
    .io_connPE_3_pop_bits(stealNW_TQ_io_connPE_3_pop_bits),
    .io_connPE_4_push_ready(stealNW_TQ_io_connPE_4_push_ready),
    .io_connPE_4_push_valid(stealNW_TQ_io_connPE_4_push_valid),
    .io_connPE_4_push_bits(stealNW_TQ_io_connPE_4_push_bits),
    .io_connPE_4_pop_ready(stealNW_TQ_io_connPE_4_pop_ready),
    .io_connPE_4_pop_valid(stealNW_TQ_io_connPE_4_pop_valid),
    .io_connPE_4_pop_bits(stealNW_TQ_io_connPE_4_pop_bits),
    .io_connPE_5_push_ready(stealNW_TQ_io_connPE_5_push_ready),
    .io_connPE_5_push_valid(stealNW_TQ_io_connPE_5_push_valid),
    .io_connPE_5_push_bits(stealNW_TQ_io_connPE_5_push_bits),
    .io_connPE_5_pop_ready(stealNW_TQ_io_connPE_5_pop_ready),
    .io_connPE_5_pop_valid(stealNW_TQ_io_connPE_5_pop_valid),
    .io_connPE_5_pop_bits(stealNW_TQ_io_connPE_5_pop_bits),
    .io_connPE_6_push_ready(stealNW_TQ_io_connPE_6_push_ready),
    .io_connPE_6_push_valid(stealNW_TQ_io_connPE_6_push_valid),
    .io_connPE_6_push_bits(stealNW_TQ_io_connPE_6_push_bits),
    .io_connPE_6_pop_ready(stealNW_TQ_io_connPE_6_pop_ready),
    .io_connPE_6_pop_valid(stealNW_TQ_io_connPE_6_pop_valid),
    .io_connPE_6_pop_bits(stealNW_TQ_io_connPE_6_pop_bits),
    .io_connPE_7_push_ready(stealNW_TQ_io_connPE_7_push_ready),
    .io_connPE_7_push_valid(stealNW_TQ_io_connPE_7_push_valid),
    .io_connPE_7_push_bits(stealNW_TQ_io_connPE_7_push_bits),
    .io_connPE_7_pop_ready(stealNW_TQ_io_connPE_7_pop_ready),
    .io_connPE_7_pop_valid(stealNW_TQ_io_connPE_7_pop_valid),
    .io_connPE_7_pop_bits(stealNW_TQ_io_connPE_7_pop_bits),
    .io_connPE_8_push_ready(stealNW_TQ_io_connPE_8_push_ready),
    .io_connPE_8_push_valid(stealNW_TQ_io_connPE_8_push_valid),
    .io_connPE_8_push_bits(stealNW_TQ_io_connPE_8_push_bits),
    .io_connPE_8_pop_ready(stealNW_TQ_io_connPE_8_pop_ready),
    .io_connPE_8_pop_valid(stealNW_TQ_io_connPE_8_pop_valid),
    .io_connPE_8_pop_bits(stealNW_TQ_io_connPE_8_pop_bits),
    .io_connPE_9_push_ready(stealNW_TQ_io_connPE_9_push_ready),
    .io_connPE_9_push_valid(stealNW_TQ_io_connPE_9_push_valid),
    .io_connPE_9_push_bits(stealNW_TQ_io_connPE_9_push_bits),
    .io_connPE_9_pop_ready(stealNW_TQ_io_connPE_9_pop_ready),
    .io_connPE_9_pop_valid(stealNW_TQ_io_connPE_9_pop_valid),
    .io_connPE_9_pop_bits(stealNW_TQ_io_connPE_9_pop_bits),
    .io_connPE_10_push_ready(stealNW_TQ_io_connPE_10_push_ready),
    .io_connPE_10_push_valid(stealNW_TQ_io_connPE_10_push_valid),
    .io_connPE_10_push_bits(stealNW_TQ_io_connPE_10_push_bits),
    .io_connPE_10_pop_ready(stealNW_TQ_io_connPE_10_pop_ready),
    .io_connPE_10_pop_valid(stealNW_TQ_io_connPE_10_pop_valid),
    .io_connPE_10_pop_bits(stealNW_TQ_io_connPE_10_pop_bits),
    .io_connPE_11_push_ready(stealNW_TQ_io_connPE_11_push_ready),
    .io_connPE_11_push_valid(stealNW_TQ_io_connPE_11_push_valid),
    .io_connPE_11_push_bits(stealNW_TQ_io_connPE_11_push_bits),
    .io_connPE_11_pop_ready(stealNW_TQ_io_connPE_11_pop_ready),
    .io_connPE_11_pop_valid(stealNW_TQ_io_connPE_11_pop_valid),
    .io_connPE_11_pop_bits(stealNW_TQ_io_connPE_11_pop_bits),
    .io_connPE_12_push_ready(stealNW_TQ_io_connPE_12_push_ready),
    .io_connPE_12_push_valid(stealNW_TQ_io_connPE_12_push_valid),
    .io_connPE_12_push_bits(stealNW_TQ_io_connPE_12_push_bits),
    .io_connPE_12_pop_ready(stealNW_TQ_io_connPE_12_pop_ready),
    .io_connPE_12_pop_valid(stealNW_TQ_io_connPE_12_pop_valid),
    .io_connPE_12_pop_bits(stealNW_TQ_io_connPE_12_pop_bits),
    .io_connPE_13_push_ready(stealNW_TQ_io_connPE_13_push_ready),
    .io_connPE_13_push_valid(stealNW_TQ_io_connPE_13_push_valid),
    .io_connPE_13_push_bits(stealNW_TQ_io_connPE_13_push_bits),
    .io_connPE_13_pop_ready(stealNW_TQ_io_connPE_13_pop_ready),
    .io_connPE_13_pop_valid(stealNW_TQ_io_connPE_13_pop_valid),
    .io_connPE_13_pop_bits(stealNW_TQ_io_connPE_13_pop_bits),
    .io_connPE_14_push_ready(stealNW_TQ_io_connPE_14_push_ready),
    .io_connPE_14_push_valid(stealNW_TQ_io_connPE_14_push_valid),
    .io_connPE_14_push_bits(stealNW_TQ_io_connPE_14_push_bits),
    .io_connPE_14_pop_ready(stealNW_TQ_io_connPE_14_pop_ready),
    .io_connPE_14_pop_valid(stealNW_TQ_io_connPE_14_pop_valid),
    .io_connPE_14_pop_bits(stealNW_TQ_io_connPE_14_pop_bits),
    .io_connPE_15_push_ready(stealNW_TQ_io_connPE_15_push_ready),
    .io_connPE_15_push_valid(stealNW_TQ_io_connPE_15_push_valid),
    .io_connPE_15_push_bits(stealNW_TQ_io_connPE_15_push_bits),
    .io_connPE_15_pop_ready(stealNW_TQ_io_connPE_15_pop_ready),
    .io_connPE_15_pop_valid(stealNW_TQ_io_connPE_15_pop_valid),
    .io_connPE_15_pop_bits(stealNW_TQ_io_connPE_15_pop_bits),
    .io_connPE_16_push_ready(stealNW_TQ_io_connPE_16_push_ready),
    .io_connPE_16_push_valid(stealNW_TQ_io_connPE_16_push_valid),
    .io_connPE_16_push_bits(stealNW_TQ_io_connPE_16_push_bits),
    .io_connPE_16_pop_ready(stealNW_TQ_io_connPE_16_pop_ready),
    .io_connPE_16_pop_valid(stealNW_TQ_io_connPE_16_pop_valid),
    .io_connPE_16_pop_bits(stealNW_TQ_io_connPE_16_pop_bits),
    .io_connPE_17_push_ready(stealNW_TQ_io_connPE_17_push_ready),
    .io_connPE_17_push_valid(stealNW_TQ_io_connPE_17_push_valid),
    .io_connPE_17_push_bits(stealNW_TQ_io_connPE_17_push_bits),
    .io_connPE_17_pop_ready(stealNW_TQ_io_connPE_17_pop_ready),
    .io_connPE_17_pop_valid(stealNW_TQ_io_connPE_17_pop_valid),
    .io_connPE_17_pop_bits(stealNW_TQ_io_connPE_17_pop_bits),
    .io_connPE_18_push_ready(stealNW_TQ_io_connPE_18_push_ready),
    .io_connPE_18_push_valid(stealNW_TQ_io_connPE_18_push_valid),
    .io_connPE_18_push_bits(stealNW_TQ_io_connPE_18_push_bits),
    .io_connPE_18_pop_ready(stealNW_TQ_io_connPE_18_pop_ready),
    .io_connPE_18_pop_valid(stealNW_TQ_io_connPE_18_pop_valid),
    .io_connPE_18_pop_bits(stealNW_TQ_io_connPE_18_pop_bits),
    .io_connPE_19_push_ready(stealNW_TQ_io_connPE_19_push_ready),
    .io_connPE_19_push_valid(stealNW_TQ_io_connPE_19_push_valid),
    .io_connPE_19_push_bits(stealNW_TQ_io_connPE_19_push_bits),
    .io_connPE_19_pop_ready(stealNW_TQ_io_connPE_19_pop_ready),
    .io_connPE_19_pop_valid(stealNW_TQ_io_connPE_19_pop_valid),
    .io_connPE_19_pop_bits(stealNW_TQ_io_connPE_19_pop_bits),
    .io_connPE_20_push_ready(stealNW_TQ_io_connPE_20_push_ready),
    .io_connPE_20_push_valid(stealNW_TQ_io_connPE_20_push_valid),
    .io_connPE_20_push_bits(stealNW_TQ_io_connPE_20_push_bits),
    .io_connPE_20_pop_ready(stealNW_TQ_io_connPE_20_pop_ready),
    .io_connPE_20_pop_valid(stealNW_TQ_io_connPE_20_pop_valid),
    .io_connPE_20_pop_bits(stealNW_TQ_io_connPE_20_pop_bits),
    .io_connPE_21_push_ready(stealNW_TQ_io_connPE_21_push_ready),
    .io_connPE_21_push_valid(stealNW_TQ_io_connPE_21_push_valid),
    .io_connPE_21_push_bits(stealNW_TQ_io_connPE_21_push_bits),
    .io_connPE_21_pop_ready(stealNW_TQ_io_connPE_21_pop_ready),
    .io_connPE_21_pop_valid(stealNW_TQ_io_connPE_21_pop_valid),
    .io_connPE_21_pop_bits(stealNW_TQ_io_connPE_21_pop_bits),
    .io_connPE_22_push_ready(stealNW_TQ_io_connPE_22_push_ready),
    .io_connPE_22_push_valid(stealNW_TQ_io_connPE_22_push_valid),
    .io_connPE_22_push_bits(stealNW_TQ_io_connPE_22_push_bits),
    .io_connPE_22_pop_ready(stealNW_TQ_io_connPE_22_pop_ready),
    .io_connPE_22_pop_valid(stealNW_TQ_io_connPE_22_pop_valid),
    .io_connPE_22_pop_bits(stealNW_TQ_io_connPE_22_pop_bits),
    .io_connPE_23_push_ready(stealNW_TQ_io_connPE_23_push_ready),
    .io_connPE_23_push_valid(stealNW_TQ_io_connPE_23_push_valid),
    .io_connPE_23_push_bits(stealNW_TQ_io_connPE_23_push_bits),
    .io_connPE_23_pop_ready(stealNW_TQ_io_connPE_23_pop_ready),
    .io_connPE_23_pop_valid(stealNW_TQ_io_connPE_23_pop_valid),
    .io_connPE_23_pop_bits(stealNW_TQ_io_connPE_23_pop_bits),
    .io_connPE_24_push_ready(stealNW_TQ_io_connPE_24_push_ready),
    .io_connPE_24_push_valid(stealNW_TQ_io_connPE_24_push_valid),
    .io_connPE_24_push_bits(stealNW_TQ_io_connPE_24_push_bits),
    .io_connPE_24_pop_ready(stealNW_TQ_io_connPE_24_pop_ready),
    .io_connPE_24_pop_valid(stealNW_TQ_io_connPE_24_pop_valid),
    .io_connPE_24_pop_bits(stealNW_TQ_io_connPE_24_pop_bits),
    .io_connPE_25_push_ready(stealNW_TQ_io_connPE_25_push_ready),
    .io_connPE_25_push_valid(stealNW_TQ_io_connPE_25_push_valid),
    .io_connPE_25_push_bits(stealNW_TQ_io_connPE_25_push_bits),
    .io_connPE_25_pop_ready(stealNW_TQ_io_connPE_25_pop_ready),
    .io_connPE_25_pop_valid(stealNW_TQ_io_connPE_25_pop_valid),
    .io_connPE_25_pop_bits(stealNW_TQ_io_connPE_25_pop_bits),
    .io_connPE_26_push_ready(stealNW_TQ_io_connPE_26_push_ready),
    .io_connPE_26_push_valid(stealNW_TQ_io_connPE_26_push_valid),
    .io_connPE_26_push_bits(stealNW_TQ_io_connPE_26_push_bits),
    .io_connPE_26_pop_ready(stealNW_TQ_io_connPE_26_pop_ready),
    .io_connPE_26_pop_valid(stealNW_TQ_io_connPE_26_pop_valid),
    .io_connPE_26_pop_bits(stealNW_TQ_io_connPE_26_pop_bits),
    .io_connPE_27_push_ready(stealNW_TQ_io_connPE_27_push_ready),
    .io_connPE_27_push_valid(stealNW_TQ_io_connPE_27_push_valid),
    .io_connPE_27_push_bits(stealNW_TQ_io_connPE_27_push_bits),
    .io_connPE_27_pop_ready(stealNW_TQ_io_connPE_27_pop_ready),
    .io_connPE_27_pop_valid(stealNW_TQ_io_connPE_27_pop_valid),
    .io_connPE_27_pop_bits(stealNW_TQ_io_connPE_27_pop_bits),
    .io_connPE_28_push_ready(stealNW_TQ_io_connPE_28_push_ready),
    .io_connPE_28_push_valid(stealNW_TQ_io_connPE_28_push_valid),
    .io_connPE_28_push_bits(stealNW_TQ_io_connPE_28_push_bits),
    .io_connPE_28_pop_ready(stealNW_TQ_io_connPE_28_pop_ready),
    .io_connPE_28_pop_valid(stealNW_TQ_io_connPE_28_pop_valid),
    .io_connPE_28_pop_bits(stealNW_TQ_io_connPE_28_pop_bits),
    .io_connPE_29_push_ready(stealNW_TQ_io_connPE_29_push_ready),
    .io_connPE_29_push_valid(stealNW_TQ_io_connPE_29_push_valid),
    .io_connPE_29_push_bits(stealNW_TQ_io_connPE_29_push_bits),
    .io_connPE_29_pop_ready(stealNW_TQ_io_connPE_29_pop_ready),
    .io_connPE_29_pop_valid(stealNW_TQ_io_connPE_29_pop_valid),
    .io_connPE_29_pop_bits(stealNW_TQ_io_connPE_29_pop_bits),
    .io_connPE_30_push_ready(stealNW_TQ_io_connPE_30_push_ready),
    .io_connPE_30_push_valid(stealNW_TQ_io_connPE_30_push_valid),
    .io_connPE_30_push_bits(stealNW_TQ_io_connPE_30_push_bits),
    .io_connPE_30_pop_ready(stealNW_TQ_io_connPE_30_pop_ready),
    .io_connPE_30_pop_valid(stealNW_TQ_io_connPE_30_pop_valid),
    .io_connPE_30_pop_bits(stealNW_TQ_io_connPE_30_pop_bits),
    .io_connPE_31_push_ready(stealNW_TQ_io_connPE_31_push_ready),
    .io_connPE_31_push_valid(stealNW_TQ_io_connPE_31_push_valid),
    .io_connPE_31_push_bits(stealNW_TQ_io_connPE_31_push_bits),
    .io_connPE_31_pop_ready(stealNW_TQ_io_connPE_31_pop_ready),
    .io_connPE_31_pop_valid(stealNW_TQ_io_connPE_31_pop_valid),
    .io_connPE_31_pop_bits(stealNW_TQ_io_connPE_31_pop_bits),
    .io_connPE_32_push_ready(stealNW_TQ_io_connPE_32_push_ready),
    .io_connPE_32_push_valid(stealNW_TQ_io_connPE_32_push_valid),
    .io_connPE_32_push_bits(stealNW_TQ_io_connPE_32_push_bits),
    .io_connPE_32_pop_ready(stealNW_TQ_io_connPE_32_pop_ready),
    .io_connPE_32_pop_valid(stealNW_TQ_io_connPE_32_pop_valid),
    .io_connPE_32_pop_bits(stealNW_TQ_io_connPE_32_pop_bits),
    .io_connPE_33_push_ready(stealNW_TQ_io_connPE_33_push_ready),
    .io_connPE_33_push_valid(stealNW_TQ_io_connPE_33_push_valid),
    .io_connPE_33_push_bits(stealNW_TQ_io_connPE_33_push_bits),
    .io_connPE_33_pop_ready(stealNW_TQ_io_connPE_33_pop_ready),
    .io_connPE_33_pop_valid(stealNW_TQ_io_connPE_33_pop_valid),
    .io_connPE_33_pop_bits(stealNW_TQ_io_connPE_33_pop_bits),
    .io_connPE_34_push_ready(stealNW_TQ_io_connPE_34_push_ready),
    .io_connPE_34_push_valid(stealNW_TQ_io_connPE_34_push_valid),
    .io_connPE_34_push_bits(stealNW_TQ_io_connPE_34_push_bits),
    .io_connPE_34_pop_ready(stealNW_TQ_io_connPE_34_pop_ready),
    .io_connPE_34_pop_valid(stealNW_TQ_io_connPE_34_pop_valid),
    .io_connPE_34_pop_bits(stealNW_TQ_io_connPE_34_pop_bits),
    .io_connPE_35_push_ready(stealNW_TQ_io_connPE_35_push_ready),
    .io_connPE_35_push_valid(stealNW_TQ_io_connPE_35_push_valid),
    .io_connPE_35_push_bits(stealNW_TQ_io_connPE_35_push_bits),
    .io_connPE_35_pop_ready(stealNW_TQ_io_connPE_35_pop_ready),
    .io_connPE_35_pop_valid(stealNW_TQ_io_connPE_35_pop_valid),
    .io_connPE_35_pop_bits(stealNW_TQ_io_connPE_35_pop_bits),
    .io_connPE_36_push_ready(stealNW_TQ_io_connPE_36_push_ready),
    .io_connPE_36_push_valid(stealNW_TQ_io_connPE_36_push_valid),
    .io_connPE_36_push_bits(stealNW_TQ_io_connPE_36_push_bits),
    .io_connPE_36_pop_ready(stealNW_TQ_io_connPE_36_pop_ready),
    .io_connPE_36_pop_valid(stealNW_TQ_io_connPE_36_pop_valid),
    .io_connPE_36_pop_bits(stealNW_TQ_io_connPE_36_pop_bits),
    .io_connPE_37_push_ready(stealNW_TQ_io_connPE_37_push_ready),
    .io_connPE_37_push_valid(stealNW_TQ_io_connPE_37_push_valid),
    .io_connPE_37_push_bits(stealNW_TQ_io_connPE_37_push_bits),
    .io_connPE_37_pop_ready(stealNW_TQ_io_connPE_37_pop_ready),
    .io_connPE_37_pop_valid(stealNW_TQ_io_connPE_37_pop_valid),
    .io_connPE_37_pop_bits(stealNW_TQ_io_connPE_37_pop_bits),
    .io_connPE_38_push_ready(stealNW_TQ_io_connPE_38_push_ready),
    .io_connPE_38_push_valid(stealNW_TQ_io_connPE_38_push_valid),
    .io_connPE_38_push_bits(stealNW_TQ_io_connPE_38_push_bits),
    .io_connPE_38_pop_ready(stealNW_TQ_io_connPE_38_pop_ready),
    .io_connPE_38_pop_valid(stealNW_TQ_io_connPE_38_pop_valid),
    .io_connPE_38_pop_bits(stealNW_TQ_io_connPE_38_pop_bits),
    .io_connPE_39_push_ready(stealNW_TQ_io_connPE_39_push_ready),
    .io_connPE_39_push_valid(stealNW_TQ_io_connPE_39_push_valid),
    .io_connPE_39_push_bits(stealNW_TQ_io_connPE_39_push_bits),
    .io_connPE_39_pop_ready(stealNW_TQ_io_connPE_39_pop_ready),
    .io_connPE_39_pop_valid(stealNW_TQ_io_connPE_39_pop_valid),
    .io_connPE_39_pop_bits(stealNW_TQ_io_connPE_39_pop_bits),
    .io_connPE_40_push_ready(stealNW_TQ_io_connPE_40_push_ready),
    .io_connPE_40_push_valid(stealNW_TQ_io_connPE_40_push_valid),
    .io_connPE_40_push_bits(stealNW_TQ_io_connPE_40_push_bits),
    .io_connPE_40_pop_ready(stealNW_TQ_io_connPE_40_pop_ready),
    .io_connPE_40_pop_valid(stealNW_TQ_io_connPE_40_pop_valid),
    .io_connPE_40_pop_bits(stealNW_TQ_io_connPE_40_pop_bits),
    .io_connPE_41_push_ready(stealNW_TQ_io_connPE_41_push_ready),
    .io_connPE_41_push_valid(stealNW_TQ_io_connPE_41_push_valid),
    .io_connPE_41_push_bits(stealNW_TQ_io_connPE_41_push_bits),
    .io_connPE_41_pop_ready(stealNW_TQ_io_connPE_41_pop_ready),
    .io_connPE_41_pop_valid(stealNW_TQ_io_connPE_41_pop_valid),
    .io_connPE_41_pop_bits(stealNW_TQ_io_connPE_41_pop_bits),
    .io_connPE_42_push_ready(stealNW_TQ_io_connPE_42_push_ready),
    .io_connPE_42_push_valid(stealNW_TQ_io_connPE_42_push_valid),
    .io_connPE_42_push_bits(stealNW_TQ_io_connPE_42_push_bits),
    .io_connPE_42_pop_ready(stealNW_TQ_io_connPE_42_pop_ready),
    .io_connPE_42_pop_valid(stealNW_TQ_io_connPE_42_pop_valid),
    .io_connPE_42_pop_bits(stealNW_TQ_io_connPE_42_pop_bits),
    .io_connPE_43_push_ready(stealNW_TQ_io_connPE_43_push_ready),
    .io_connPE_43_push_valid(stealNW_TQ_io_connPE_43_push_valid),
    .io_connPE_43_push_bits(stealNW_TQ_io_connPE_43_push_bits),
    .io_connPE_43_pop_ready(stealNW_TQ_io_connPE_43_pop_ready),
    .io_connPE_43_pop_valid(stealNW_TQ_io_connPE_43_pop_valid),
    .io_connPE_43_pop_bits(stealNW_TQ_io_connPE_43_pop_bits),
    .io_connPE_44_push_ready(stealNW_TQ_io_connPE_44_push_ready),
    .io_connPE_44_push_valid(stealNW_TQ_io_connPE_44_push_valid),
    .io_connPE_44_push_bits(stealNW_TQ_io_connPE_44_push_bits),
    .io_connPE_44_pop_ready(stealNW_TQ_io_connPE_44_pop_ready),
    .io_connPE_44_pop_valid(stealNW_TQ_io_connPE_44_pop_valid),
    .io_connPE_44_pop_bits(stealNW_TQ_io_connPE_44_pop_bits),
    .io_connPE_45_push_ready(stealNW_TQ_io_connPE_45_push_ready),
    .io_connPE_45_push_valid(stealNW_TQ_io_connPE_45_push_valid),
    .io_connPE_45_push_bits(stealNW_TQ_io_connPE_45_push_bits),
    .io_connPE_45_pop_ready(stealNW_TQ_io_connPE_45_pop_ready),
    .io_connPE_45_pop_valid(stealNW_TQ_io_connPE_45_pop_valid),
    .io_connPE_45_pop_bits(stealNW_TQ_io_connPE_45_pop_bits),
    .io_connPE_46_push_ready(stealNW_TQ_io_connPE_46_push_ready),
    .io_connPE_46_push_valid(stealNW_TQ_io_connPE_46_push_valid),
    .io_connPE_46_push_bits(stealNW_TQ_io_connPE_46_push_bits),
    .io_connPE_46_pop_ready(stealNW_TQ_io_connPE_46_pop_ready),
    .io_connPE_46_pop_valid(stealNW_TQ_io_connPE_46_pop_valid),
    .io_connPE_46_pop_bits(stealNW_TQ_io_connPE_46_pop_bits),
    .io_connPE_47_push_ready(stealNW_TQ_io_connPE_47_push_ready),
    .io_connPE_47_push_valid(stealNW_TQ_io_connPE_47_push_valid),
    .io_connPE_47_push_bits(stealNW_TQ_io_connPE_47_push_bits),
    .io_connPE_47_pop_ready(stealNW_TQ_io_connPE_47_pop_ready),
    .io_connPE_47_pop_valid(stealNW_TQ_io_connPE_47_pop_valid),
    .io_connPE_47_pop_bits(stealNW_TQ_io_connPE_47_pop_bits),
    .io_connPE_48_push_ready(stealNW_TQ_io_connPE_48_push_ready),
    .io_connPE_48_push_valid(stealNW_TQ_io_connPE_48_push_valid),
    .io_connPE_48_push_bits(stealNW_TQ_io_connPE_48_push_bits),
    .io_connPE_48_pop_ready(stealNW_TQ_io_connPE_48_pop_ready),
    .io_connPE_48_pop_valid(stealNW_TQ_io_connPE_48_pop_valid),
    .io_connPE_48_pop_bits(stealNW_TQ_io_connPE_48_pop_bits),
    .io_connPE_49_push_ready(stealNW_TQ_io_connPE_49_push_ready),
    .io_connPE_49_push_valid(stealNW_TQ_io_connPE_49_push_valid),
    .io_connPE_49_push_bits(stealNW_TQ_io_connPE_49_push_bits),
    .io_connPE_49_pop_ready(stealNW_TQ_io_connPE_49_pop_ready),
    .io_connPE_49_pop_valid(stealNW_TQ_io_connPE_49_pop_valid),
    .io_connPE_49_pop_bits(stealNW_TQ_io_connPE_49_pop_bits),
    .io_connPE_50_push_ready(stealNW_TQ_io_connPE_50_push_ready),
    .io_connPE_50_push_valid(stealNW_TQ_io_connPE_50_push_valid),
    .io_connPE_50_push_bits(stealNW_TQ_io_connPE_50_push_bits),
    .io_connPE_50_pop_ready(stealNW_TQ_io_connPE_50_pop_ready),
    .io_connPE_50_pop_valid(stealNW_TQ_io_connPE_50_pop_valid),
    .io_connPE_50_pop_bits(stealNW_TQ_io_connPE_50_pop_bits),
    .io_connPE_51_push_ready(stealNW_TQ_io_connPE_51_push_ready),
    .io_connPE_51_push_valid(stealNW_TQ_io_connPE_51_push_valid),
    .io_connPE_51_push_bits(stealNW_TQ_io_connPE_51_push_bits),
    .io_connPE_51_pop_ready(stealNW_TQ_io_connPE_51_pop_ready),
    .io_connPE_51_pop_valid(stealNW_TQ_io_connPE_51_pop_valid),
    .io_connPE_51_pop_bits(stealNW_TQ_io_connPE_51_pop_bits),
    .io_connPE_52_push_ready(stealNW_TQ_io_connPE_52_push_ready),
    .io_connPE_52_push_valid(stealNW_TQ_io_connPE_52_push_valid),
    .io_connPE_52_push_bits(stealNW_TQ_io_connPE_52_push_bits),
    .io_connPE_52_pop_ready(stealNW_TQ_io_connPE_52_pop_ready),
    .io_connPE_52_pop_valid(stealNW_TQ_io_connPE_52_pop_valid),
    .io_connPE_52_pop_bits(stealNW_TQ_io_connPE_52_pop_bits),
    .io_connPE_53_push_ready(stealNW_TQ_io_connPE_53_push_ready),
    .io_connPE_53_push_valid(stealNW_TQ_io_connPE_53_push_valid),
    .io_connPE_53_push_bits(stealNW_TQ_io_connPE_53_push_bits),
    .io_connPE_53_pop_ready(stealNW_TQ_io_connPE_53_pop_ready),
    .io_connPE_53_pop_valid(stealNW_TQ_io_connPE_53_pop_valid),
    .io_connPE_53_pop_bits(stealNW_TQ_io_connPE_53_pop_bits),
    .io_connPE_54_push_ready(stealNW_TQ_io_connPE_54_push_ready),
    .io_connPE_54_push_valid(stealNW_TQ_io_connPE_54_push_valid),
    .io_connPE_54_push_bits(stealNW_TQ_io_connPE_54_push_bits),
    .io_connPE_54_pop_ready(stealNW_TQ_io_connPE_54_pop_ready),
    .io_connPE_54_pop_valid(stealNW_TQ_io_connPE_54_pop_valid),
    .io_connPE_54_pop_bits(stealNW_TQ_io_connPE_54_pop_bits),
    .io_connPE_55_push_ready(stealNW_TQ_io_connPE_55_push_ready),
    .io_connPE_55_push_valid(stealNW_TQ_io_connPE_55_push_valid),
    .io_connPE_55_push_bits(stealNW_TQ_io_connPE_55_push_bits),
    .io_connPE_55_pop_ready(stealNW_TQ_io_connPE_55_pop_ready),
    .io_connPE_55_pop_valid(stealNW_TQ_io_connPE_55_pop_valid),
    .io_connPE_55_pop_bits(stealNW_TQ_io_connPE_55_pop_bits),
    .io_connPE_56_push_ready(stealNW_TQ_io_connPE_56_push_ready),
    .io_connPE_56_push_valid(stealNW_TQ_io_connPE_56_push_valid),
    .io_connPE_56_push_bits(stealNW_TQ_io_connPE_56_push_bits),
    .io_connPE_56_pop_ready(stealNW_TQ_io_connPE_56_pop_ready),
    .io_connPE_56_pop_valid(stealNW_TQ_io_connPE_56_pop_valid),
    .io_connPE_56_pop_bits(stealNW_TQ_io_connPE_56_pop_bits),
    .io_connPE_57_push_ready(stealNW_TQ_io_connPE_57_push_ready),
    .io_connPE_57_push_valid(stealNW_TQ_io_connPE_57_push_valid),
    .io_connPE_57_push_bits(stealNW_TQ_io_connPE_57_push_bits),
    .io_connPE_57_pop_ready(stealNW_TQ_io_connPE_57_pop_ready),
    .io_connPE_57_pop_valid(stealNW_TQ_io_connPE_57_pop_valid),
    .io_connPE_57_pop_bits(stealNW_TQ_io_connPE_57_pop_bits),
    .io_connPE_58_push_ready(stealNW_TQ_io_connPE_58_push_ready),
    .io_connPE_58_push_valid(stealNW_TQ_io_connPE_58_push_valid),
    .io_connPE_58_push_bits(stealNW_TQ_io_connPE_58_push_bits),
    .io_connPE_58_pop_ready(stealNW_TQ_io_connPE_58_pop_ready),
    .io_connPE_58_pop_valid(stealNW_TQ_io_connPE_58_pop_valid),
    .io_connPE_58_pop_bits(stealNW_TQ_io_connPE_58_pop_bits),
    .io_connPE_59_push_ready(stealNW_TQ_io_connPE_59_push_ready),
    .io_connPE_59_push_valid(stealNW_TQ_io_connPE_59_push_valid),
    .io_connPE_59_push_bits(stealNW_TQ_io_connPE_59_push_bits),
    .io_connPE_59_pop_ready(stealNW_TQ_io_connPE_59_pop_ready),
    .io_connPE_59_pop_valid(stealNW_TQ_io_connPE_59_pop_valid),
    .io_connPE_59_pop_bits(stealNW_TQ_io_connPE_59_pop_bits),
    .io_connPE_60_push_ready(stealNW_TQ_io_connPE_60_push_ready),
    .io_connPE_60_push_valid(stealNW_TQ_io_connPE_60_push_valid),
    .io_connPE_60_push_bits(stealNW_TQ_io_connPE_60_push_bits),
    .io_connPE_60_pop_ready(stealNW_TQ_io_connPE_60_pop_ready),
    .io_connPE_60_pop_valid(stealNW_TQ_io_connPE_60_pop_valid),
    .io_connPE_60_pop_bits(stealNW_TQ_io_connPE_60_pop_bits),
    .io_connPE_61_push_ready(stealNW_TQ_io_connPE_61_push_ready),
    .io_connPE_61_push_valid(stealNW_TQ_io_connPE_61_push_valid),
    .io_connPE_61_push_bits(stealNW_TQ_io_connPE_61_push_bits),
    .io_connPE_61_pop_ready(stealNW_TQ_io_connPE_61_pop_ready),
    .io_connPE_61_pop_valid(stealNW_TQ_io_connPE_61_pop_valid),
    .io_connPE_61_pop_bits(stealNW_TQ_io_connPE_61_pop_bits),
    .io_connPE_62_push_ready(stealNW_TQ_io_connPE_62_push_ready),
    .io_connPE_62_push_valid(stealNW_TQ_io_connPE_62_push_valid),
    .io_connPE_62_push_bits(stealNW_TQ_io_connPE_62_push_bits),
    .io_connPE_62_pop_ready(stealNW_TQ_io_connPE_62_pop_ready),
    .io_connPE_62_pop_valid(stealNW_TQ_io_connPE_62_pop_valid),
    .io_connPE_62_pop_bits(stealNW_TQ_io_connPE_62_pop_bits),
    .io_connPE_63_push_ready(stealNW_TQ_io_connPE_63_push_ready),
    .io_connPE_63_push_valid(stealNW_TQ_io_connPE_63_push_valid),
    .io_connPE_63_push_bits(stealNW_TQ_io_connPE_63_push_bits),
    .io_connPE_63_pop_ready(stealNW_TQ_io_connPE_63_pop_ready),
    .io_connPE_63_pop_valid(stealNW_TQ_io_connPE_63_pop_valid),
    .io_connPE_63_pop_bits(stealNW_TQ_io_connPE_63_pop_bits),
    .io_connVSS_0_ctrl_serveStealReq_ready(stealNW_TQ_io_connVSS_0_ctrl_serveStealReq_ready),
    .io_connVSS_0_ctrl_serveStealReq_valid(stealNW_TQ_io_connVSS_0_ctrl_serveStealReq_valid),
    .io_connVSS_0_data_availableTask_ready(stealNW_TQ_io_connVSS_0_data_availableTask_ready),
    .io_connVSS_0_data_availableTask_valid(stealNW_TQ_io_connVSS_0_data_availableTask_valid),
    .io_connVSS_0_data_availableTask_bits(stealNW_TQ_io_connVSS_0_data_availableTask_bits),
    .io_connVSS_0_data_qOutTask_ready(stealNW_TQ_io_connVSS_0_data_qOutTask_ready),
    .io_connVSS_0_data_qOutTask_valid(stealNW_TQ_io_connVSS_0_data_qOutTask_valid),
    .io_connVSS_0_data_qOutTask_bits(stealNW_TQ_io_connVSS_0_data_qOutTask_bits),
    .io_connVAS_0_ctrl_serveStealReq_ready(stealNW_TQ_io_connVAS_0_ctrl_serveStealReq_ready),
    .io_connVAS_0_ctrl_serveStealReq_valid(stealNW_TQ_io_connVAS_0_ctrl_serveStealReq_valid),
    .io_connVAS_0_data_qOutTask_ready(stealNW_TQ_io_connVAS_0_data_qOutTask_ready),
    .io_connVAS_0_data_qOutTask_valid(stealNW_TQ_io_connVAS_0_data_qOutTask_valid),
    .io_connVAS_0_data_qOutTask_bits(stealNW_TQ_io_connVAS_0_data_qOutTask_bits),
    .io_connVAS_1_ctrl_serveStealReq_ready(stealNW_TQ_io_connVAS_1_ctrl_serveStealReq_ready),
    .io_connVAS_1_ctrl_serveStealReq_valid(stealNW_TQ_io_connVAS_1_ctrl_serveStealReq_valid),
    .io_connVAS_1_data_qOutTask_ready(stealNW_TQ_io_connVAS_1_data_qOutTask_ready),
    .io_connVAS_1_data_qOutTask_valid(stealNW_TQ_io_connVAS_1_data_qOutTask_valid),
    .io_connVAS_1_data_qOutTask_bits(stealNW_TQ_io_connVAS_1_data_qOutTask_bits),
    .io_ntwDataUnitOccupancyVSS_0(stealNW_TQ_io_ntwDataUnitOccupancyVSS_0)
  );
  virtualStealServer virtualStealServers_0 ( // @[stealSide.scala 66:75]
    .clock(virtualStealServers_0_clock),
    .reset(virtualStealServers_0_reset),
    .io_connNetwork_ctrl_serveStealReq_ready(virtualStealServers_0_io_connNetwork_ctrl_serveStealReq_ready),
    .io_connNetwork_ctrl_serveStealReq_valid(virtualStealServers_0_io_connNetwork_ctrl_serveStealReq_valid),
    .io_connNetwork_data_availableTask_ready(virtualStealServers_0_io_connNetwork_data_availableTask_ready),
    .io_connNetwork_data_availableTask_valid(virtualStealServers_0_io_connNetwork_data_availableTask_valid),
    .io_connNetwork_data_availableTask_bits(virtualStealServers_0_io_connNetwork_data_availableTask_bits),
    .io_connNetwork_data_qOutTask_ready(virtualStealServers_0_io_connNetwork_data_qOutTask_ready),
    .io_connNetwork_data_qOutTask_valid(virtualStealServers_0_io_connNetwork_data_qOutTask_valid),
    .io_connNetwork_data_qOutTask_bits(virtualStealServers_0_io_connNetwork_data_qOutTask_bits),
    .io_axi_mgmt_ARREADY(virtualStealServers_0_io_axi_mgmt_ARREADY),
    .io_axi_mgmt_ARVALID(virtualStealServers_0_io_axi_mgmt_ARVALID),
    .io_axi_mgmt_ARADDR(virtualStealServers_0_io_axi_mgmt_ARADDR),
    .io_axi_mgmt_RREADY(virtualStealServers_0_io_axi_mgmt_RREADY),
    .io_axi_mgmt_RVALID(virtualStealServers_0_io_axi_mgmt_RVALID),
    .io_axi_mgmt_RDATA(virtualStealServers_0_io_axi_mgmt_RDATA),
    .io_axi_mgmt_AWREADY(virtualStealServers_0_io_axi_mgmt_AWREADY),
    .io_axi_mgmt_AWVALID(virtualStealServers_0_io_axi_mgmt_AWVALID),
    .io_axi_mgmt_AWADDR(virtualStealServers_0_io_axi_mgmt_AWADDR),
    .io_axi_mgmt_WREADY(virtualStealServers_0_io_axi_mgmt_WREADY),
    .io_axi_mgmt_WVALID(virtualStealServers_0_io_axi_mgmt_WVALID),
    .io_axi_mgmt_WDATA(virtualStealServers_0_io_axi_mgmt_WDATA),
    .io_axi_mgmt_WSTRB(virtualStealServers_0_io_axi_mgmt_WSTRB),
    .io_axi_mgmt_BREADY(virtualStealServers_0_io_axi_mgmt_BREADY),
    .io_axi_mgmt_BVALID(virtualStealServers_0_io_axi_mgmt_BVALID),
    .io_read_address_ready(virtualStealServers_0_io_read_address_ready),
    .io_read_address_valid(virtualStealServers_0_io_read_address_valid),
    .io_read_address_bits(virtualStealServers_0_io_read_address_bits),
    .io_read_data_ready(virtualStealServers_0_io_read_data_ready),
    .io_read_data_valid(virtualStealServers_0_io_read_data_valid),
    .io_read_data_bits(virtualStealServers_0_io_read_data_bits),
    .io_read_burst_len(virtualStealServers_0_io_read_burst_len),
    .io_write_address_ready(virtualStealServers_0_io_write_address_ready),
    .io_write_address_valid(virtualStealServers_0_io_write_address_valid),
    .io_write_address_bits(virtualStealServers_0_io_write_address_bits),
    .io_write_data_ready(virtualStealServers_0_io_write_data_ready),
    .io_write_data_valid(virtualStealServers_0_io_write_data_valid),
    .io_write_data_bits(virtualStealServers_0_io_write_data_bits),
    .io_write_burst_len(virtualStealServers_0_io_write_burst_len),
    .io_write_last(virtualStealServers_0_io_write_last),
    .io_ntwDataUnitOccupancy(virtualStealServers_0_io_ntwDataUnitOccupancy)
  );
  readyValidMem vssRvm_0 ( // @[stealSide.scala 91:68]
    .clock(vssRvm_0_clock),
    .reset(vssRvm_0_reset),
    .io_read_address_ready(vssRvm_0_io_read_address_ready),
    .io_read_address_valid(vssRvm_0_io_read_address_valid),
    .io_read_address_bits(vssRvm_0_io_read_address_bits),
    .io_read_data_ready(vssRvm_0_io_read_data_ready),
    .io_read_data_valid(vssRvm_0_io_read_data_valid),
    .io_read_data_bits(vssRvm_0_io_read_data_bits),
    .io_write_address_ready(vssRvm_0_io_write_address_ready),
    .io_write_address_valid(vssRvm_0_io_write_address_valid),
    .io_write_address_bits(vssRvm_0_io_write_address_bits),
    .io_write_data_ready(vssRvm_0_io_write_data_ready),
    .io_write_data_valid(vssRvm_0_io_write_data_valid),
    .io_write_data_bits(vssRvm_0_io_write_data_bits),
    .io_writeBurst_len(vssRvm_0_io_writeBurst_len),
    .io_writeBurst_last(vssRvm_0_io_writeBurst_last),
    .io_readBurst_len(vssRvm_0_io_readBurst_len),
    .axi_ARREADY(vssRvm_0_axi_ARREADY),
    .axi_ARVALID(vssRvm_0_axi_ARVALID),
    .axi_ARADDR(vssRvm_0_axi_ARADDR),
    .axi_ARLEN(vssRvm_0_axi_ARLEN),
    .axi_RREADY(vssRvm_0_axi_RREADY),
    .axi_RVALID(vssRvm_0_axi_RVALID),
    .axi_RDATA(vssRvm_0_axi_RDATA),
    .axi_AWREADY(vssRvm_0_axi_AWREADY),
    .axi_AWVALID(vssRvm_0_axi_AWVALID),
    .axi_AWADDR(vssRvm_0_axi_AWADDR),
    .axi_AWLEN(vssRvm_0_axi_AWLEN),
    .axi_WREADY(vssRvm_0_axi_WREADY),
    .axi_WVALID(vssRvm_0_axi_WVALID),
    .axi_WDATA(vssRvm_0_axi_WDATA),
    .axi_WLAST(vssRvm_0_axi_WLAST),
    .axi_BVALID(vssRvm_0_axi_BVALID)
  );
  assign io_axi_mgmt_vss_0_ARREADY = virtualStealServers_0_io_axi_mgmt_ARREADY; // @[stealSide.scala 87:28]
  assign io_axi_mgmt_vss_0_RVALID = virtualStealServers_0_io_axi_mgmt_RVALID; // @[stealSide.scala 87:28]
  assign io_axi_mgmt_vss_0_RDATA = virtualStealServers_0_io_axi_mgmt_RDATA; // @[stealSide.scala 87:28]
  assign io_axi_mgmt_vss_0_AWREADY = virtualStealServers_0_io_axi_mgmt_AWREADY; // @[stealSide.scala 87:28]
  assign io_axi_mgmt_vss_0_WREADY = virtualStealServers_0_io_axi_mgmt_WREADY; // @[stealSide.scala 87:28]
  assign io_axi_mgmt_vss_0_BVALID = virtualStealServers_0_io_axi_mgmt_BVALID; // @[stealSide.scala 87:28]
  assign io_vss_axi_full_0_ARVALID = vssRvm_0_axi_ARVALID; // @[stealSide.scala 102:47]
  assign io_vss_axi_full_0_ARADDR = vssRvm_0_axi_ARADDR; // @[stealSide.scala 102:47]
  assign io_vss_axi_full_0_ARLEN = vssRvm_0_axi_ARLEN; // @[stealSide.scala 102:47]
  assign io_vss_axi_full_0_RREADY = vssRvm_0_axi_RREADY; // @[stealSide.scala 102:47]
  assign io_vss_axi_full_0_AWVALID = vssRvm_0_axi_AWVALID; // @[stealSide.scala 102:47]
  assign io_vss_axi_full_0_AWADDR = vssRvm_0_axi_AWADDR; // @[stealSide.scala 102:47]
  assign io_vss_axi_full_0_AWLEN = vssRvm_0_axi_AWLEN; // @[stealSide.scala 102:47]
  assign io_vss_axi_full_0_WVALID = vssRvm_0_axi_WVALID; // @[stealSide.scala 102:47]
  assign io_vss_axi_full_0_WDATA = vssRvm_0_axi_WDATA; // @[stealSide.scala 102:47]
  assign io_vss_axi_full_0_WLAST = vssRvm_0_axi_WLAST; // @[stealSide.scala 102:47]
  assign io_taskOut_0_TVALID = stealNW_TQ_io_connPE_0_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_0_TDATA = stealNW_TQ_io_connPE_0_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_1_TVALID = stealNW_TQ_io_connPE_1_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_1_TDATA = stealNW_TQ_io_connPE_1_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_2_TVALID = stealNW_TQ_io_connPE_2_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_2_TDATA = stealNW_TQ_io_connPE_2_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_3_TVALID = stealNW_TQ_io_connPE_3_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_3_TDATA = stealNW_TQ_io_connPE_3_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_4_TVALID = stealNW_TQ_io_connPE_4_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_4_TDATA = stealNW_TQ_io_connPE_4_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_5_TVALID = stealNW_TQ_io_connPE_5_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_5_TDATA = stealNW_TQ_io_connPE_5_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_6_TVALID = stealNW_TQ_io_connPE_6_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_6_TDATA = stealNW_TQ_io_connPE_6_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_7_TVALID = stealNW_TQ_io_connPE_7_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_7_TDATA = stealNW_TQ_io_connPE_7_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_8_TVALID = stealNW_TQ_io_connPE_8_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_8_TDATA = stealNW_TQ_io_connPE_8_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_9_TVALID = stealNW_TQ_io_connPE_9_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_9_TDATA = stealNW_TQ_io_connPE_9_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_10_TVALID = stealNW_TQ_io_connPE_10_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_10_TDATA = stealNW_TQ_io_connPE_10_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_11_TVALID = stealNW_TQ_io_connPE_11_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_11_TDATA = stealNW_TQ_io_connPE_11_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_12_TVALID = stealNW_TQ_io_connPE_12_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_12_TDATA = stealNW_TQ_io_connPE_12_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_13_TVALID = stealNW_TQ_io_connPE_13_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_13_TDATA = stealNW_TQ_io_connPE_13_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_14_TVALID = stealNW_TQ_io_connPE_14_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_14_TDATA = stealNW_TQ_io_connPE_14_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_15_TVALID = stealNW_TQ_io_connPE_15_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_15_TDATA = stealNW_TQ_io_connPE_15_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_16_TVALID = stealNW_TQ_io_connPE_16_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_16_TDATA = stealNW_TQ_io_connPE_16_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_17_TVALID = stealNW_TQ_io_connPE_17_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_17_TDATA = stealNW_TQ_io_connPE_17_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_18_TVALID = stealNW_TQ_io_connPE_18_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_18_TDATA = stealNW_TQ_io_connPE_18_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_19_TVALID = stealNW_TQ_io_connPE_19_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_19_TDATA = stealNW_TQ_io_connPE_19_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_20_TVALID = stealNW_TQ_io_connPE_20_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_20_TDATA = stealNW_TQ_io_connPE_20_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_21_TVALID = stealNW_TQ_io_connPE_21_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_21_TDATA = stealNW_TQ_io_connPE_21_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_22_TVALID = stealNW_TQ_io_connPE_22_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_22_TDATA = stealNW_TQ_io_connPE_22_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_23_TVALID = stealNW_TQ_io_connPE_23_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_23_TDATA = stealNW_TQ_io_connPE_23_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_24_TVALID = stealNW_TQ_io_connPE_24_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_24_TDATA = stealNW_TQ_io_connPE_24_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_25_TVALID = stealNW_TQ_io_connPE_25_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_25_TDATA = stealNW_TQ_io_connPE_25_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_26_TVALID = stealNW_TQ_io_connPE_26_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_26_TDATA = stealNW_TQ_io_connPE_26_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_27_TVALID = stealNW_TQ_io_connPE_27_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_27_TDATA = stealNW_TQ_io_connPE_27_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_28_TVALID = stealNW_TQ_io_connPE_28_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_28_TDATA = stealNW_TQ_io_connPE_28_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_29_TVALID = stealNW_TQ_io_connPE_29_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_29_TDATA = stealNW_TQ_io_connPE_29_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_30_TVALID = stealNW_TQ_io_connPE_30_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_30_TDATA = stealNW_TQ_io_connPE_30_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_31_TVALID = stealNW_TQ_io_connPE_31_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_31_TDATA = stealNW_TQ_io_connPE_31_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_32_TVALID = stealNW_TQ_io_connPE_32_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_32_TDATA = stealNW_TQ_io_connPE_32_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_33_TVALID = stealNW_TQ_io_connPE_33_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_33_TDATA = stealNW_TQ_io_connPE_33_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_34_TVALID = stealNW_TQ_io_connPE_34_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_34_TDATA = stealNW_TQ_io_connPE_34_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_35_TVALID = stealNW_TQ_io_connPE_35_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_35_TDATA = stealNW_TQ_io_connPE_35_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_36_TVALID = stealNW_TQ_io_connPE_36_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_36_TDATA = stealNW_TQ_io_connPE_36_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_37_TVALID = stealNW_TQ_io_connPE_37_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_37_TDATA = stealNW_TQ_io_connPE_37_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_38_TVALID = stealNW_TQ_io_connPE_38_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_38_TDATA = stealNW_TQ_io_connPE_38_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_39_TVALID = stealNW_TQ_io_connPE_39_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_39_TDATA = stealNW_TQ_io_connPE_39_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_40_TVALID = stealNW_TQ_io_connPE_40_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_40_TDATA = stealNW_TQ_io_connPE_40_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_41_TVALID = stealNW_TQ_io_connPE_41_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_41_TDATA = stealNW_TQ_io_connPE_41_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_42_TVALID = stealNW_TQ_io_connPE_42_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_42_TDATA = stealNW_TQ_io_connPE_42_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_43_TVALID = stealNW_TQ_io_connPE_43_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_43_TDATA = stealNW_TQ_io_connPE_43_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_44_TVALID = stealNW_TQ_io_connPE_44_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_44_TDATA = stealNW_TQ_io_connPE_44_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_45_TVALID = stealNW_TQ_io_connPE_45_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_45_TDATA = stealNW_TQ_io_connPE_45_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_46_TVALID = stealNW_TQ_io_connPE_46_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_46_TDATA = stealNW_TQ_io_connPE_46_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_47_TVALID = stealNW_TQ_io_connPE_47_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_47_TDATA = stealNW_TQ_io_connPE_47_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_48_TVALID = stealNW_TQ_io_connPE_48_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_48_TDATA = stealNW_TQ_io_connPE_48_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_49_TVALID = stealNW_TQ_io_connPE_49_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_49_TDATA = stealNW_TQ_io_connPE_49_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_50_TVALID = stealNW_TQ_io_connPE_50_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_50_TDATA = stealNW_TQ_io_connPE_50_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_51_TVALID = stealNW_TQ_io_connPE_51_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_51_TDATA = stealNW_TQ_io_connPE_51_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_52_TVALID = stealNW_TQ_io_connPE_52_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_52_TDATA = stealNW_TQ_io_connPE_52_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_53_TVALID = stealNW_TQ_io_connPE_53_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_53_TDATA = stealNW_TQ_io_connPE_53_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_54_TVALID = stealNW_TQ_io_connPE_54_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_54_TDATA = stealNW_TQ_io_connPE_54_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_55_TVALID = stealNW_TQ_io_connPE_55_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_55_TDATA = stealNW_TQ_io_connPE_55_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_56_TVALID = stealNW_TQ_io_connPE_56_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_56_TDATA = stealNW_TQ_io_connPE_56_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_57_TVALID = stealNW_TQ_io_connPE_57_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_57_TDATA = stealNW_TQ_io_connPE_57_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_58_TVALID = stealNW_TQ_io_connPE_58_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_58_TDATA = stealNW_TQ_io_connPE_58_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_59_TVALID = stealNW_TQ_io_connPE_59_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_59_TDATA = stealNW_TQ_io_connPE_59_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_60_TVALID = stealNW_TQ_io_connPE_60_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_60_TDATA = stealNW_TQ_io_connPE_60_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_61_TVALID = stealNW_TQ_io_connPE_61_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_61_TDATA = stealNW_TQ_io_connPE_61_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_62_TVALID = stealNW_TQ_io_connPE_62_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_62_TDATA = stealNW_TQ_io_connPE_62_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskOut_63_TVALID = stealNW_TQ_io_connPE_63_pop_valid; // @[stealSide.scala 107:39]
  assign io_taskOut_63_TDATA = stealNW_TQ_io_connPE_63_pop_bits; // @[stealSide.scala 107:39]
  assign io_taskIn_0_TREADY = stealNW_TQ_io_connPE_0_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_1_TREADY = stealNW_TQ_io_connPE_1_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_2_TREADY = stealNW_TQ_io_connPE_2_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_3_TREADY = stealNW_TQ_io_connPE_3_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_4_TREADY = stealNW_TQ_io_connPE_4_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_5_TREADY = stealNW_TQ_io_connPE_5_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_6_TREADY = stealNW_TQ_io_connPE_6_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_7_TREADY = stealNW_TQ_io_connPE_7_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_8_TREADY = stealNW_TQ_io_connPE_8_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_9_TREADY = stealNW_TQ_io_connPE_9_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_10_TREADY = stealNW_TQ_io_connPE_10_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_11_TREADY = stealNW_TQ_io_connPE_11_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_12_TREADY = stealNW_TQ_io_connPE_12_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_13_TREADY = stealNW_TQ_io_connPE_13_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_14_TREADY = stealNW_TQ_io_connPE_14_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_15_TREADY = stealNW_TQ_io_connPE_15_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_16_TREADY = stealNW_TQ_io_connPE_16_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_17_TREADY = stealNW_TQ_io_connPE_17_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_18_TREADY = stealNW_TQ_io_connPE_18_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_19_TREADY = stealNW_TQ_io_connPE_19_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_20_TREADY = stealNW_TQ_io_connPE_20_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_21_TREADY = stealNW_TQ_io_connPE_21_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_22_TREADY = stealNW_TQ_io_connPE_22_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_23_TREADY = stealNW_TQ_io_connPE_23_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_24_TREADY = stealNW_TQ_io_connPE_24_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_25_TREADY = stealNW_TQ_io_connPE_25_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_26_TREADY = stealNW_TQ_io_connPE_26_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_27_TREADY = stealNW_TQ_io_connPE_27_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_28_TREADY = stealNW_TQ_io_connPE_28_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_29_TREADY = stealNW_TQ_io_connPE_29_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_30_TREADY = stealNW_TQ_io_connPE_30_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_31_TREADY = stealNW_TQ_io_connPE_31_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_32_TREADY = stealNW_TQ_io_connPE_32_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_33_TREADY = stealNW_TQ_io_connPE_33_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_34_TREADY = stealNW_TQ_io_connPE_34_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_35_TREADY = stealNW_TQ_io_connPE_35_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_36_TREADY = stealNW_TQ_io_connPE_36_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_37_TREADY = stealNW_TQ_io_connPE_37_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_38_TREADY = stealNW_TQ_io_connPE_38_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_39_TREADY = stealNW_TQ_io_connPE_39_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_40_TREADY = stealNW_TQ_io_connPE_40_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_41_TREADY = stealNW_TQ_io_connPE_41_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_42_TREADY = stealNW_TQ_io_connPE_42_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_43_TREADY = stealNW_TQ_io_connPE_43_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_44_TREADY = stealNW_TQ_io_connPE_44_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_45_TREADY = stealNW_TQ_io_connPE_45_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_46_TREADY = stealNW_TQ_io_connPE_46_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_47_TREADY = stealNW_TQ_io_connPE_47_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_48_TREADY = stealNW_TQ_io_connPE_48_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_49_TREADY = stealNW_TQ_io_connPE_49_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_50_TREADY = stealNW_TQ_io_connPE_50_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_51_TREADY = stealNW_TQ_io_connPE_51_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_52_TREADY = stealNW_TQ_io_connPE_52_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_53_TREADY = stealNW_TQ_io_connPE_53_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_54_TREADY = stealNW_TQ_io_connPE_54_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_55_TREADY = stealNW_TQ_io_connPE_55_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_56_TREADY = stealNW_TQ_io_connPE_56_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_57_TREADY = stealNW_TQ_io_connPE_57_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_58_TREADY = stealNW_TQ_io_connPE_58_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_59_TREADY = stealNW_TQ_io_connPE_59_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_60_TREADY = stealNW_TQ_io_connPE_60_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_61_TREADY = stealNW_TQ_io_connPE_61_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_62_TREADY = stealNW_TQ_io_connPE_62_push_ready; // @[stealSide.scala 109:43]
  assign io_taskIn_63_TREADY = stealNW_TQ_io_connPE_63_push_ready; // @[stealSide.scala 109:43]
  assign connSyncSide_0_ctrl_serveStealReq_ready = stealNW_TQ_io_connVAS_0_ctrl_serveStealReq_ready; // @[stealSide.scala 118:38]
  assign connSyncSide_0_data_qOutTask_ready = stealNW_TQ_io_connVAS_0_data_qOutTask_ready; // @[stealSide.scala 118:38]
  assign connSyncSide_1_ctrl_serveStealReq_ready = stealNW_TQ_io_connVAS_1_ctrl_serveStealReq_ready; // @[stealSide.scala 118:38]
  assign connSyncSide_1_data_qOutTask_ready = stealNW_TQ_io_connVAS_1_data_qOutTask_ready; // @[stealSide.scala 118:38]
  assign stealNW_TQ_clock = clock;
  assign stealNW_TQ_reset = reset;
  assign stealNW_TQ_io_connPE_0_push_valid = io_taskIn_0_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_0_push_bits = io_taskIn_0_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_0_pop_ready = io_taskOut_0_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_1_push_valid = io_taskIn_1_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_1_push_bits = io_taskIn_1_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_1_pop_ready = io_taskOut_1_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_2_push_valid = io_taskIn_2_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_2_push_bits = io_taskIn_2_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_2_pop_ready = io_taskOut_2_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_3_push_valid = io_taskIn_3_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_3_push_bits = io_taskIn_3_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_3_pop_ready = io_taskOut_3_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_4_push_valid = io_taskIn_4_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_4_push_bits = io_taskIn_4_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_4_pop_ready = io_taskOut_4_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_5_push_valid = io_taskIn_5_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_5_push_bits = io_taskIn_5_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_5_pop_ready = io_taskOut_5_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_6_push_valid = io_taskIn_6_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_6_push_bits = io_taskIn_6_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_6_pop_ready = io_taskOut_6_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_7_push_valid = io_taskIn_7_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_7_push_bits = io_taskIn_7_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_7_pop_ready = io_taskOut_7_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_8_push_valid = io_taskIn_8_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_8_push_bits = io_taskIn_8_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_8_pop_ready = io_taskOut_8_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_9_push_valid = io_taskIn_9_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_9_push_bits = io_taskIn_9_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_9_pop_ready = io_taskOut_9_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_10_push_valid = io_taskIn_10_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_10_push_bits = io_taskIn_10_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_10_pop_ready = io_taskOut_10_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_11_push_valid = io_taskIn_11_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_11_push_bits = io_taskIn_11_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_11_pop_ready = io_taskOut_11_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_12_push_valid = io_taskIn_12_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_12_push_bits = io_taskIn_12_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_12_pop_ready = io_taskOut_12_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_13_push_valid = io_taskIn_13_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_13_push_bits = io_taskIn_13_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_13_pop_ready = io_taskOut_13_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_14_push_valid = io_taskIn_14_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_14_push_bits = io_taskIn_14_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_14_pop_ready = io_taskOut_14_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_15_push_valid = io_taskIn_15_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_15_push_bits = io_taskIn_15_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_15_pop_ready = io_taskOut_15_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_16_push_valid = io_taskIn_16_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_16_push_bits = io_taskIn_16_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_16_pop_ready = io_taskOut_16_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_17_push_valid = io_taskIn_17_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_17_push_bits = io_taskIn_17_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_17_pop_ready = io_taskOut_17_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_18_push_valid = io_taskIn_18_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_18_push_bits = io_taskIn_18_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_18_pop_ready = io_taskOut_18_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_19_push_valid = io_taskIn_19_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_19_push_bits = io_taskIn_19_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_19_pop_ready = io_taskOut_19_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_20_push_valid = io_taskIn_20_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_20_push_bits = io_taskIn_20_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_20_pop_ready = io_taskOut_20_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_21_push_valid = io_taskIn_21_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_21_push_bits = io_taskIn_21_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_21_pop_ready = io_taskOut_21_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_22_push_valid = io_taskIn_22_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_22_push_bits = io_taskIn_22_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_22_pop_ready = io_taskOut_22_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_23_push_valid = io_taskIn_23_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_23_push_bits = io_taskIn_23_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_23_pop_ready = io_taskOut_23_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_24_push_valid = io_taskIn_24_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_24_push_bits = io_taskIn_24_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_24_pop_ready = io_taskOut_24_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_25_push_valid = io_taskIn_25_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_25_push_bits = io_taskIn_25_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_25_pop_ready = io_taskOut_25_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_26_push_valid = io_taskIn_26_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_26_push_bits = io_taskIn_26_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_26_pop_ready = io_taskOut_26_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_27_push_valid = io_taskIn_27_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_27_push_bits = io_taskIn_27_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_27_pop_ready = io_taskOut_27_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_28_push_valid = io_taskIn_28_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_28_push_bits = io_taskIn_28_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_28_pop_ready = io_taskOut_28_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_29_push_valid = io_taskIn_29_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_29_push_bits = io_taskIn_29_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_29_pop_ready = io_taskOut_29_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_30_push_valid = io_taskIn_30_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_30_push_bits = io_taskIn_30_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_30_pop_ready = io_taskOut_30_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_31_push_valid = io_taskIn_31_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_31_push_bits = io_taskIn_31_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_31_pop_ready = io_taskOut_31_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_32_push_valid = io_taskIn_32_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_32_push_bits = io_taskIn_32_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_32_pop_ready = io_taskOut_32_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_33_push_valid = io_taskIn_33_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_33_push_bits = io_taskIn_33_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_33_pop_ready = io_taskOut_33_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_34_push_valid = io_taskIn_34_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_34_push_bits = io_taskIn_34_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_34_pop_ready = io_taskOut_34_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_35_push_valid = io_taskIn_35_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_35_push_bits = io_taskIn_35_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_35_pop_ready = io_taskOut_35_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_36_push_valid = io_taskIn_36_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_36_push_bits = io_taskIn_36_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_36_pop_ready = io_taskOut_36_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_37_push_valid = io_taskIn_37_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_37_push_bits = io_taskIn_37_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_37_pop_ready = io_taskOut_37_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_38_push_valid = io_taskIn_38_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_38_push_bits = io_taskIn_38_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_38_pop_ready = io_taskOut_38_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_39_push_valid = io_taskIn_39_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_39_push_bits = io_taskIn_39_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_39_pop_ready = io_taskOut_39_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_40_push_valid = io_taskIn_40_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_40_push_bits = io_taskIn_40_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_40_pop_ready = io_taskOut_40_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_41_push_valid = io_taskIn_41_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_41_push_bits = io_taskIn_41_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_41_pop_ready = io_taskOut_41_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_42_push_valid = io_taskIn_42_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_42_push_bits = io_taskIn_42_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_42_pop_ready = io_taskOut_42_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_43_push_valid = io_taskIn_43_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_43_push_bits = io_taskIn_43_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_43_pop_ready = io_taskOut_43_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_44_push_valid = io_taskIn_44_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_44_push_bits = io_taskIn_44_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_44_pop_ready = io_taskOut_44_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_45_push_valid = io_taskIn_45_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_45_push_bits = io_taskIn_45_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_45_pop_ready = io_taskOut_45_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_46_push_valid = io_taskIn_46_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_46_push_bits = io_taskIn_46_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_46_pop_ready = io_taskOut_46_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_47_push_valid = io_taskIn_47_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_47_push_bits = io_taskIn_47_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_47_pop_ready = io_taskOut_47_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_48_push_valid = io_taskIn_48_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_48_push_bits = io_taskIn_48_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_48_pop_ready = io_taskOut_48_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_49_push_valid = io_taskIn_49_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_49_push_bits = io_taskIn_49_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_49_pop_ready = io_taskOut_49_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_50_push_valid = io_taskIn_50_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_50_push_bits = io_taskIn_50_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_50_pop_ready = io_taskOut_50_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_51_push_valid = io_taskIn_51_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_51_push_bits = io_taskIn_51_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_51_pop_ready = io_taskOut_51_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_52_push_valid = io_taskIn_52_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_52_push_bits = io_taskIn_52_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_52_pop_ready = io_taskOut_52_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_53_push_valid = io_taskIn_53_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_53_push_bits = io_taskIn_53_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_53_pop_ready = io_taskOut_53_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_54_push_valid = io_taskIn_54_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_54_push_bits = io_taskIn_54_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_54_pop_ready = io_taskOut_54_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_55_push_valid = io_taskIn_55_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_55_push_bits = io_taskIn_55_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_55_pop_ready = io_taskOut_55_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_56_push_valid = io_taskIn_56_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_56_push_bits = io_taskIn_56_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_56_pop_ready = io_taskOut_56_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_57_push_valid = io_taskIn_57_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_57_push_bits = io_taskIn_57_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_57_pop_ready = io_taskOut_57_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_58_push_valid = io_taskIn_58_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_58_push_bits = io_taskIn_58_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_58_pop_ready = io_taskOut_58_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_59_push_valid = io_taskIn_59_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_59_push_bits = io_taskIn_59_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_59_pop_ready = io_taskOut_59_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_60_push_valid = io_taskIn_60_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_60_push_bits = io_taskIn_60_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_60_pop_ready = io_taskOut_60_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_61_push_valid = io_taskIn_61_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_61_push_bits = io_taskIn_61_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_61_pop_ready = io_taskOut_61_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_62_push_valid = io_taskIn_62_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_62_push_bits = io_taskIn_62_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_62_pop_ready = io_taskOut_62_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connPE_63_push_valid = io_taskIn_63_TVALID; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_63_push_bits = io_taskIn_63_TDATA; // @[stealSide.scala 109:43]
  assign stealNW_TQ_io_connPE_63_pop_ready = io_taskOut_63_TREADY; // @[stealSide.scala 107:39]
  assign stealNW_TQ_io_connVSS_0_ctrl_serveStealReq_valid =
    virtualStealServers_0_io_connNetwork_ctrl_serveStealReq_valid; // @[stealSide.scala 103:47]
  assign stealNW_TQ_io_connVSS_0_data_availableTask_ready =
    virtualStealServers_0_io_connNetwork_data_availableTask_ready; // @[stealSide.scala 103:47]
  assign stealNW_TQ_io_connVSS_0_data_qOutTask_valid = virtualStealServers_0_io_connNetwork_data_qOutTask_valid; // @[stealSide.scala 103:47]
  assign stealNW_TQ_io_connVSS_0_data_qOutTask_bits = virtualStealServers_0_io_connNetwork_data_qOutTask_bits; // @[stealSide.scala 103:47]
  assign stealNW_TQ_io_connVAS_0_ctrl_serveStealReq_valid = connSyncSide_0_ctrl_serveStealReq_valid; // @[stealSide.scala 118:38]
  assign stealNW_TQ_io_connVAS_0_data_qOutTask_valid = connSyncSide_0_data_qOutTask_valid; // @[stealSide.scala 118:38]
  assign stealNW_TQ_io_connVAS_0_data_qOutTask_bits = connSyncSide_0_data_qOutTask_bits; // @[stealSide.scala 118:38]
  assign stealNW_TQ_io_connVAS_1_ctrl_serveStealReq_valid = connSyncSide_1_ctrl_serveStealReq_valid; // @[stealSide.scala 118:38]
  assign stealNW_TQ_io_connVAS_1_data_qOutTask_valid = connSyncSide_1_data_qOutTask_valid; // @[stealSide.scala 118:38]
  assign stealNW_TQ_io_connVAS_1_data_qOutTask_bits = connSyncSide_1_data_qOutTask_bits; // @[stealSide.scala 118:38]
  assign virtualStealServers_0_clock = clock;
  assign virtualStealServers_0_reset = reset;
  assign virtualStealServers_0_io_connNetwork_ctrl_serveStealReq_ready =
    stealNW_TQ_io_connVSS_0_ctrl_serveStealReq_ready; // @[stealSide.scala 103:47]
  assign virtualStealServers_0_io_connNetwork_data_availableTask_valid =
    stealNW_TQ_io_connVSS_0_data_availableTask_valid; // @[stealSide.scala 103:47]
  assign virtualStealServers_0_io_connNetwork_data_availableTask_bits = stealNW_TQ_io_connVSS_0_data_availableTask_bits; // @[stealSide.scala 103:47]
  assign virtualStealServers_0_io_connNetwork_data_qOutTask_ready = stealNW_TQ_io_connVSS_0_data_qOutTask_ready; // @[stealSide.scala 103:47]
  assign virtualStealServers_0_io_axi_mgmt_ARVALID = io_axi_mgmt_vss_0_ARVALID; // @[stealSide.scala 87:28]
  assign virtualStealServers_0_io_axi_mgmt_ARADDR = io_axi_mgmt_vss_0_ARADDR; // @[stealSide.scala 87:28]
  assign virtualStealServers_0_io_axi_mgmt_RREADY = io_axi_mgmt_vss_0_RREADY; // @[stealSide.scala 87:28]
  assign virtualStealServers_0_io_axi_mgmt_AWVALID = io_axi_mgmt_vss_0_AWVALID; // @[stealSide.scala 87:28]
  assign virtualStealServers_0_io_axi_mgmt_AWADDR = io_axi_mgmt_vss_0_AWADDR; // @[stealSide.scala 87:28]
  assign virtualStealServers_0_io_axi_mgmt_WVALID = io_axi_mgmt_vss_0_WVALID; // @[stealSide.scala 87:28]
  assign virtualStealServers_0_io_axi_mgmt_WDATA = io_axi_mgmt_vss_0_WDATA; // @[stealSide.scala 87:28]
  assign virtualStealServers_0_io_axi_mgmt_WSTRB = io_axi_mgmt_vss_0_WSTRB; // @[stealSide.scala 87:28]
  assign virtualStealServers_0_io_axi_mgmt_BREADY = io_axi_mgmt_vss_0_BREADY; // @[stealSide.scala 87:28]
  assign virtualStealServers_0_io_read_address_ready = vssRvm_0_io_read_address_ready; // @[stealSide.scala 95:47]
  assign virtualStealServers_0_io_read_data_valid = vssRvm_0_io_read_data_valid; // @[stealSide.scala 96:47]
  assign virtualStealServers_0_io_read_data_bits = vssRvm_0_io_read_data_bits; // @[stealSide.scala 96:47]
  assign virtualStealServers_0_io_write_address_ready = vssRvm_0_io_write_address_ready; // @[stealSide.scala 97:47]
  assign virtualStealServers_0_io_write_data_ready = vssRvm_0_io_write_data_ready; // @[stealSide.scala 98:47]
  assign virtualStealServers_0_io_ntwDataUnitOccupancy = stealNW_TQ_io_ntwDataUnitOccupancyVSS_0; // @[stealSide.scala 88:56]
  assign vssRvm_0_clock = clock;
  assign vssRvm_0_reset = reset;
  assign vssRvm_0_io_read_address_valid = virtualStealServers_0_io_read_address_valid; // @[stealSide.scala 95:47]
  assign vssRvm_0_io_read_address_bits = virtualStealServers_0_io_read_address_bits; // @[stealSide.scala 95:47]
  assign vssRvm_0_io_read_data_ready = virtualStealServers_0_io_read_data_ready; // @[stealSide.scala 96:47]
  assign vssRvm_0_io_write_address_valid = virtualStealServers_0_io_write_address_valid; // @[stealSide.scala 97:47]
  assign vssRvm_0_io_write_address_bits = virtualStealServers_0_io_write_address_bits; // @[stealSide.scala 97:47]
  assign vssRvm_0_io_write_data_valid = virtualStealServers_0_io_write_data_valid; // @[stealSide.scala 98:47]
  assign vssRvm_0_io_write_data_bits = virtualStealServers_0_io_write_data_bits; // @[stealSide.scala 98:47]
  assign vssRvm_0_io_writeBurst_len = virtualStealServers_0_io_write_burst_len; // @[stealSide.scala 100:47]
  assign vssRvm_0_io_writeBurst_last = virtualStealServers_0_io_write_last; // @[stealSide.scala 101:47]
  assign vssRvm_0_io_readBurst_len = virtualStealServers_0_io_read_burst_len; // @[stealSide.scala 99:47]
  assign vssRvm_0_axi_ARREADY = io_vss_axi_full_0_ARREADY; // @[stealSide.scala 102:47]
  assign vssRvm_0_axi_RVALID = io_vss_axi_full_0_RVALID; // @[stealSide.scala 102:47]
  assign vssRvm_0_axi_RDATA = io_vss_axi_full_0_RDATA; // @[stealSide.scala 102:47]
  assign vssRvm_0_axi_AWREADY = io_vss_axi_full_0_AWREADY; // @[stealSide.scala 102:47]
  assign vssRvm_0_axi_WREADY = io_vss_axi_full_0_WREADY; // @[stealSide.scala 102:47]
  assign vssRvm_0_axi_BVALID = io_vss_axi_full_0_BVALID; // @[stealSide.scala 102:47]
endmodule
module contAddrNtwUnitCAS(
  input         clock,
  input         reset,
  output        io_addressIn1_ready,
  input         io_addressIn1_valid,
  input  [63:0] io_addressIn1_bits,
  input         io_addressOut_ready,
  output        io_addressOut_valid,
  output [63:0] io_addressOut_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] stateReg; // @[contAddrNtwUnitCAS.scala 24:30]
  reg [63:0] addressReg; // @[contAddrNtwUnitCAS.scala 25:30]
  reg  priorityReg; // @[contAddrNtwUnitCAS.scala 26:30]
  wire  _T = stateReg == 2'h0; // @[contAddrNtwUnitCAS.scala 34:19]
  wire  _priorityReg_T = ~priorityReg; // @[contAddrNtwUnitCAS.scala 38:28]
  wire  _GEN_0 = io_addressIn1_valid ? _priorityReg_T : priorityReg; // @[contAddrNtwUnitCAS.scala 42:40 44:25 26:30]
  wire  _T_1 = stateReg == 2'h1; // @[contAddrNtwUnitCAS.scala 49:25]
  wire  _T_2 = stateReg == 2'h2; // @[contAddrNtwUnitCAS.scala 64:25]
  wire  _GEN_10 = priorityReg ? 1'h0 : 1'h1; // @[contAddrNtwUnitCAS.scala 68:30 70:26 74:26]
  wire [1:0] _GEN_11 = io_addressOut_ready ? {{1'd0}, _GEN_10} : stateReg; // @[contAddrNtwUnitCAS.scala 24:30 66:35]
  wire  _GEN_13 = stateReg == 2'h1 ? _GEN_0 : priorityReg; // @[contAddrNtwUnitCAS.scala 26:30 49:51]
  wire  _GEN_16 = stateReg == 2'h0 ? _GEN_0 : _GEN_13; // @[contAddrNtwUnitCAS.scala 34:44]
  wire  _GEN_21 = _T_1 ? 1'h0 : _T_2; // @[contAddrNtwUnitCAS.scala 30:28 86:50]
  assign io_addressIn1_ready = _T ? 1'h0 : _T_1; // @[contAddrNtwUnitCAS.scala 29:29 82:44]
  assign io_addressOut_valid = _T ? 1'h0 : _GEN_21; // @[contAddrNtwUnitCAS.scala 30:28 82:44]
  assign io_addressOut_bits = addressReg; // @[contAddrNtwUnitCAS.scala 31:28]
  always @(posedge clock) begin
    if (reset) begin // @[contAddrNtwUnitCAS.scala 24:30]
      stateReg <= 2'h0; // @[contAddrNtwUnitCAS.scala 24:30]
    end else if (stateReg == 2'h0) begin // @[contAddrNtwUnitCAS.scala 34:44]
      if (io_addressIn1_valid) begin // @[contAddrNtwUnitCAS.scala 42:40]
        stateReg <= 2'h1; // @[contAddrNtwUnitCAS.scala 45:25]
      end
    end else if (stateReg == 2'h1) begin // @[contAddrNtwUnitCAS.scala 49:51]
      if (io_addressIn1_valid) begin // @[contAddrNtwUnitCAS.scala 51:34]
        stateReg <= 2'h2; // @[contAddrNtwUnitCAS.scala 54:25]
      end
    end else if (stateReg == 2'h2) begin // @[contAddrNtwUnitCAS.scala 64:44]
      stateReg <= _GEN_11;
    end
    if (reset) begin // @[contAddrNtwUnitCAS.scala 25:30]
      addressReg <= 64'h0; // @[contAddrNtwUnitCAS.scala 25:30]
    end else if (!(stateReg == 2'h0)) begin // @[contAddrNtwUnitCAS.scala 34:44]
      if (stateReg == 2'h1) begin // @[contAddrNtwUnitCAS.scala 49:51]
        if (io_addressIn1_valid) begin // @[contAddrNtwUnitCAS.scala 51:34]
          addressReg <= io_addressIn1_bits; // @[contAddrNtwUnitCAS.scala 55:25]
        end
      end
    end
    priorityReg <= reset | _GEN_16; // @[contAddrNtwUnitCAS.scala 26:{30,30}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  addressReg = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  priorityReg = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module contAddrNtwUnit(
  input         clock,
  input         reset,
  output        io_addressIn_ready,
  input         io_addressIn_valid,
  input  [63:0] io_addressIn_bits,
  input         io_addressOut_ready,
  output        io_addressOut_valid,
  output [63:0] io_addressOut_bits,
  input         io_casAddressOut_ready,
  output        io_casAddressOut_valid,
  output [63:0] io_casAddressOut_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  stateReg; // @[contAddrNtwUnit.scala 22:30]
  reg [63:0] addressReg; // @[contAddrNtwUnit.scala 23:30]
  reg  priorityReg; // @[contAddrNtwUnit.scala 24:30]
  wire  _T = ~stateReg; // @[contAddrNtwUnit.scala 33:19]
  wire  _GEN_1 = io_addressIn_valid | stateReg; // @[contAddrNtwUnit.scala 34:33 36:24 22:30]
  wire  _GEN_2 = io_addressOut_ready | io_casAddressOut_ready ? 1'h0 : stateReg; // @[contAddrNtwUnit.scala 39:60 40:22 22:30]
  wire  _GEN_3 = io_addressOut_ready | io_casAddressOut_ready ? ~priorityReg : priorityReg; // @[contAddrNtwUnit.scala 39:60 41:25 24:30]
  wire  _GEN_4 = stateReg & _GEN_2; // @[contAddrNtwUnit.scala 38:44 44:18]
  wire  _GEN_5 = stateReg ? _GEN_3 : priorityReg; // @[contAddrNtwUnit.scala 24:30 38:44]
  wire  _GEN_8 = ~stateReg ? priorityReg : _GEN_5; // @[contAddrNtwUnit.scala 24:30 33:43]
  wire  _GEN_11 = priorityReg & io_casAddressOut_ready; // @[contAddrNtwUnit.scala 29:28 51:30]
  wire  _GEN_12 = priorityReg ? 1'h0 : io_addressOut_ready; // @[contAddrNtwUnit.scala 27:28 51:30]
  wire  _GEN_13 = io_casAddressOut_ready ? 1'h0 : io_addressOut_ready; // @[contAddrNtwUnit.scala 27:28 61:41]
  wire  _GEN_14 = io_addressOut_ready & io_casAddressOut_ready ? _GEN_11 : io_casAddressOut_ready; // @[contAddrNtwUnit.scala 50:60]
  wire  _GEN_15 = io_addressOut_ready & io_casAddressOut_ready ? _GEN_12 : _GEN_13; // @[contAddrNtwUnit.scala 50:60]
  wire  _GEN_16 = stateReg & _GEN_14; // @[contAddrNtwUnit.scala 29:28 49:44]
  wire  _GEN_17 = stateReg & _GEN_15; // @[contAddrNtwUnit.scala 27:28 49:44]
  assign io_addressIn_ready = ~stateReg; // @[contAddrNtwUnit.scala 47:19]
  assign io_addressOut_valid = _T ? 1'h0 : _GEN_17; // @[contAddrNtwUnit.scala 27:28 47:43]
  assign io_addressOut_bits = addressReg; // @[contAddrNtwUnit.scala 28:28]
  assign io_casAddressOut_valid = _T ? 1'h0 : _GEN_16; // @[contAddrNtwUnit.scala 29:28 47:43]
  assign io_casAddressOut_bits = addressReg; // @[contAddrNtwUnit.scala 30:28]
  always @(posedge clock) begin
    if (reset) begin // @[contAddrNtwUnit.scala 22:30]
      stateReg <= 1'h0; // @[contAddrNtwUnit.scala 22:30]
    end else if (~stateReg) begin // @[contAddrNtwUnit.scala 33:43]
      stateReg <= _GEN_1;
    end else begin
      stateReg <= _GEN_4;
    end
    if (reset) begin // @[contAddrNtwUnit.scala 23:30]
      addressReg <= 64'h0; // @[contAddrNtwUnit.scala 23:30]
    end else if (~stateReg) begin // @[contAddrNtwUnit.scala 33:43]
      if (io_addressIn_valid) begin // @[contAddrNtwUnit.scala 34:33]
        addressReg <= io_addressIn_bits; // @[contAddrNtwUnit.scala 35:24]
      end
    end
    priorityReg <= reset | _GEN_8; // @[contAddrNtwUnit.scala 24:{30,30}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  addressReg = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  priorityReg = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module contAddrServer(
  input         clock,
  input         reset,
  output        io_addressIn_ready,
  input         io_addressIn_valid,
  input  [63:0] io_addressIn_bits,
  input         io_addressOut_ready,
  output        io_addressOut_valid,
  output [63:0] io_addressOut_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  stateReg; // @[contAddrServer.scala 21:27]
  reg [63:0] addressReg; // @[contAddrServer.scala 22:29]
  wire  _T = ~stateReg; // @[contAddrServer.scala 28:19]
  wire  _GEN_0 = io_addressIn_valid | stateReg; // @[contAddrServer.scala 29:33 30:24 21:27]
  wire  _GEN_2 = io_addressOut_ready ? 1'h0 : stateReg; // @[contAddrServer.scala 34:34 35:24 21:27]
  wire  _GEN_3 = stateReg & _GEN_2; // @[contAddrServer.scala 33:53 38:18]
  assign io_addressIn_ready = ~stateReg; // @[contAddrServer.scala 41:19]
  assign io_addressOut_valid = _T ? 1'h0 : stateReg; // @[contAddrServer.scala 25:25 41:43]
  assign io_addressOut_bits = addressReg; // @[contAddrServer.scala 24:25]
  always @(posedge clock) begin
    if (reset) begin // @[contAddrServer.scala 21:27]
      stateReg <= 1'h0; // @[contAddrServer.scala 21:27]
    end else if (~stateReg) begin // @[contAddrServer.scala 28:43]
      stateReg <= _GEN_0;
    end else begin
      stateReg <= _GEN_3;
    end
    if (reset) begin // @[contAddrServer.scala 22:29]
      addressReg <= 64'h0; // @[contAddrServer.scala 22:29]
    end else if (~stateReg) begin // @[contAddrServer.scala 28:43]
      if (io_addressIn_valid) begin // @[contAddrServer.scala 29:33]
        addressReg <= io_addressIn_bits; // @[contAddrServer.scala 31:24]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  addressReg = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_4(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram [0:7]; // @[Decoupled.scala 275:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 275:95]
  wire [2:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 275:95]
  wire [63:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 275:95]
  wire [63:0] ram_MPORT_data; // @[Decoupled.scala 275:95]
  wire [2:0] ram_MPORT_addr; // @[Decoupled.scala 275:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 275:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 275:95]
  reg [2:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [2:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 278:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 279:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 280:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 281:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 52:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 52:35]
  wire [2:0] _value_T_1 = enq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  wire [2:0] _value_T_3 = deq_ptr_value + 3'h1; // @[Counter.scala 77:24]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 275:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 305:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 304:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 312:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 275:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 288:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 3'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 292:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 278:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 278:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 295:27]
      maybe_full <= do_enq; // @[Decoupled.scala 296:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module contQueue(
  input         clock,
  input         reset,
  output        io_addressIn_ready,
  input         io_addressIn_valid,
  input  [63:0] io_addressIn_bits,
  input         io_addressOut_ready,
  output        io_addressOut_valid,
  output [63:0] io_addressOut_bits
);
  wire  q_clock; // @[contQueue.scala 13:19]
  wire  q_reset; // @[contQueue.scala 13:19]
  wire  q_io_enq_ready; // @[contQueue.scala 13:19]
  wire  q_io_enq_valid; // @[contQueue.scala 13:19]
  wire [63:0] q_io_enq_bits; // @[contQueue.scala 13:19]
  wire  q_io_deq_ready; // @[contQueue.scala 13:19]
  wire  q_io_deq_valid; // @[contQueue.scala 13:19]
  wire [63:0] q_io_deq_bits; // @[contQueue.scala 13:19]
  Queue_4 q ( // @[contQueue.scala 13:19]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits(q_io_enq_bits),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits(q_io_deq_bits)
  );
  assign io_addressIn_ready = q_io_enq_ready; // @[contQueue.scala 15:14]
  assign io_addressOut_valid = q_io_deq_valid; // @[contQueue.scala 16:19]
  assign io_addressOut_bits = q_io_deq_bits; // @[contQueue.scala 16:19]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_addressIn_valid; // @[contQueue.scala 15:14]
  assign q_io_enq_bits = io_addressIn_bits; // @[contQueue.scala 15:14]
  assign q_io_deq_ready = io_addressOut_ready; // @[contQueue.scala 16:19]
endmodule
module contNetwork(
  input         clock,
  input         reset,
  output        io_connVCAS_0_ready,
  input         io_connVCAS_0_valid,
  input  [63:0] io_connVCAS_0_bits,
  input         io_connPE_0_ready,
  output        io_connPE_0_valid,
  output [63:0] io_connPE_0_bits,
  input         io_connPE_1_ready,
  output        io_connPE_1_valid,
  output [63:0] io_connPE_1_bits,
  input         io_connPE_2_ready,
  output        io_connPE_2_valid,
  output [63:0] io_connPE_2_bits,
  input         io_connPE_3_ready,
  output        io_connPE_3_valid,
  output [63:0] io_connPE_3_bits,
  input         io_connPE_4_ready,
  output        io_connPE_4_valid,
  output [63:0] io_connPE_4_bits,
  input         io_connPE_5_ready,
  output        io_connPE_5_valid,
  output [63:0] io_connPE_5_bits,
  input         io_connPE_6_ready,
  output        io_connPE_6_valid,
  output [63:0] io_connPE_6_bits,
  input         io_connPE_7_ready,
  output        io_connPE_7_valid,
  output [63:0] io_connPE_7_bits,
  input         io_connPE_8_ready,
  output        io_connPE_8_valid,
  output [63:0] io_connPE_8_bits,
  input         io_connPE_9_ready,
  output        io_connPE_9_valid,
  output [63:0] io_connPE_9_bits,
  input         io_connPE_10_ready,
  output        io_connPE_10_valid,
  output [63:0] io_connPE_10_bits,
  input         io_connPE_11_ready,
  output        io_connPE_11_valid,
  output [63:0] io_connPE_11_bits,
  input         io_connPE_12_ready,
  output        io_connPE_12_valid,
  output [63:0] io_connPE_12_bits,
  input         io_connPE_13_ready,
  output        io_connPE_13_valid,
  output [63:0] io_connPE_13_bits,
  input         io_connPE_14_ready,
  output        io_connPE_14_valid,
  output [63:0] io_connPE_14_bits,
  input         io_connPE_15_ready,
  output        io_connPE_15_valid,
  output [63:0] io_connPE_15_bits,
  input         io_connPE_16_ready,
  output        io_connPE_16_valid,
  output [63:0] io_connPE_16_bits,
  input         io_connPE_17_ready,
  output        io_connPE_17_valid,
  output [63:0] io_connPE_17_bits,
  input         io_connPE_18_ready,
  output        io_connPE_18_valid,
  output [63:0] io_connPE_18_bits,
  input         io_connPE_19_ready,
  output        io_connPE_19_valid,
  output [63:0] io_connPE_19_bits,
  input         io_connPE_20_ready,
  output        io_connPE_20_valid,
  output [63:0] io_connPE_20_bits,
  input         io_connPE_21_ready,
  output        io_connPE_21_valid,
  output [63:0] io_connPE_21_bits,
  input         io_connPE_22_ready,
  output        io_connPE_22_valid,
  output [63:0] io_connPE_22_bits,
  input         io_connPE_23_ready,
  output        io_connPE_23_valid,
  output [63:0] io_connPE_23_bits,
  input         io_connPE_24_ready,
  output        io_connPE_24_valid,
  output [63:0] io_connPE_24_bits,
  input         io_connPE_25_ready,
  output        io_connPE_25_valid,
  output [63:0] io_connPE_25_bits,
  input         io_connPE_26_ready,
  output        io_connPE_26_valid,
  output [63:0] io_connPE_26_bits,
  input         io_connPE_27_ready,
  output        io_connPE_27_valid,
  output [63:0] io_connPE_27_bits,
  input         io_connPE_28_ready,
  output        io_connPE_28_valid,
  output [63:0] io_connPE_28_bits,
  input         io_connPE_29_ready,
  output        io_connPE_29_valid,
  output [63:0] io_connPE_29_bits,
  input         io_connPE_30_ready,
  output        io_connPE_30_valid,
  output [63:0] io_connPE_30_bits,
  input         io_connPE_31_ready,
  output        io_connPE_31_valid,
  output [63:0] io_connPE_31_bits,
  input         io_connPE_32_ready,
  output        io_connPE_32_valid,
  output [63:0] io_connPE_32_bits,
  input         io_connPE_33_ready,
  output        io_connPE_33_valid,
  output [63:0] io_connPE_33_bits,
  input         io_connPE_34_ready,
  output        io_connPE_34_valid,
  output [63:0] io_connPE_34_bits,
  input         io_connPE_35_ready,
  output        io_connPE_35_valid,
  output [63:0] io_connPE_35_bits,
  input         io_connPE_36_ready,
  output        io_connPE_36_valid,
  output [63:0] io_connPE_36_bits,
  input         io_connPE_37_ready,
  output        io_connPE_37_valid,
  output [63:0] io_connPE_37_bits,
  input         io_connPE_38_ready,
  output        io_connPE_38_valid,
  output [63:0] io_connPE_38_bits,
  input         io_connPE_39_ready,
  output        io_connPE_39_valid,
  output [63:0] io_connPE_39_bits,
  input         io_connPE_40_ready,
  output        io_connPE_40_valid,
  output [63:0] io_connPE_40_bits,
  input         io_connPE_41_ready,
  output        io_connPE_41_valid,
  output [63:0] io_connPE_41_bits,
  input         io_connPE_42_ready,
  output        io_connPE_42_valid,
  output [63:0] io_connPE_42_bits,
  input         io_connPE_43_ready,
  output        io_connPE_43_valid,
  output [63:0] io_connPE_43_bits,
  input         io_connPE_44_ready,
  output        io_connPE_44_valid,
  output [63:0] io_connPE_44_bits,
  input         io_connPE_45_ready,
  output        io_connPE_45_valid,
  output [63:0] io_connPE_45_bits,
  input         io_connPE_46_ready,
  output        io_connPE_46_valid,
  output [63:0] io_connPE_46_bits,
  input         io_connPE_47_ready,
  output        io_connPE_47_valid,
  output [63:0] io_connPE_47_bits,
  input         io_connPE_48_ready,
  output        io_connPE_48_valid,
  output [63:0] io_connPE_48_bits,
  input         io_connPE_49_ready,
  output        io_connPE_49_valid,
  output [63:0] io_connPE_49_bits,
  input         io_connPE_50_ready,
  output        io_connPE_50_valid,
  output [63:0] io_connPE_50_bits,
  input         io_connPE_51_ready,
  output        io_connPE_51_valid,
  output [63:0] io_connPE_51_bits,
  input         io_connPE_52_ready,
  output        io_connPE_52_valid,
  output [63:0] io_connPE_52_bits,
  input         io_connPE_53_ready,
  output        io_connPE_53_valid,
  output [63:0] io_connPE_53_bits,
  input         io_connPE_54_ready,
  output        io_connPE_54_valid,
  output [63:0] io_connPE_54_bits,
  input         io_connPE_55_ready,
  output        io_connPE_55_valid,
  output [63:0] io_connPE_55_bits,
  input         io_connPE_56_ready,
  output        io_connPE_56_valid,
  output [63:0] io_connPE_56_bits,
  input         io_connPE_57_ready,
  output        io_connPE_57_valid,
  output [63:0] io_connPE_57_bits,
  input         io_connPE_58_ready,
  output        io_connPE_58_valid,
  output [63:0] io_connPE_58_bits,
  input         io_connPE_59_ready,
  output        io_connPE_59_valid,
  output [63:0] io_connPE_59_bits,
  input         io_connPE_60_ready,
  output        io_connPE_60_valid,
  output [63:0] io_connPE_60_bits,
  input         io_connPE_61_ready,
  output        io_connPE_61_valid,
  output [63:0] io_connPE_61_bits,
  input         io_connPE_62_ready,
  output        io_connPE_62_valid,
  output [63:0] io_connPE_62_bits,
  input         io_connPE_63_ready,
  output        io_connPE_63_valid,
  output [63:0] io_connPE_63_bits
);
  wire  vcasNetworkUnits_0_clock; // @[contNetwork.scala 15:55]
  wire  vcasNetworkUnits_0_reset; // @[contNetwork.scala 15:55]
  wire  vcasNetworkUnits_0_io_addressIn1_ready; // @[contNetwork.scala 15:55]
  wire  vcasNetworkUnits_0_io_addressIn1_valid; // @[contNetwork.scala 15:55]
  wire [63:0] vcasNetworkUnits_0_io_addressIn1_bits; // @[contNetwork.scala 15:55]
  wire  vcasNetworkUnits_0_io_addressOut_ready; // @[contNetwork.scala 15:55]
  wire  vcasNetworkUnits_0_io_addressOut_valid; // @[contNetwork.scala 15:55]
  wire [63:0] vcasNetworkUnits_0_io_addressOut_bits; // @[contNetwork.scala 15:55]
  wire  networkUnits_0_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_0_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_0_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_0_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_0_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_0_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_0_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_0_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_0_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_0_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_0_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_1_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_1_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_1_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_1_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_1_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_1_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_1_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_1_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_1_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_1_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_1_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_2_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_2_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_2_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_2_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_2_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_2_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_2_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_2_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_2_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_2_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_2_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_3_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_3_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_3_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_3_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_3_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_3_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_3_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_3_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_3_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_3_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_3_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_4_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_4_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_4_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_4_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_4_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_4_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_4_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_4_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_4_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_4_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_4_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_5_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_5_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_5_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_5_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_5_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_5_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_5_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_5_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_5_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_5_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_5_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_6_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_6_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_6_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_6_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_6_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_6_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_6_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_6_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_6_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_6_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_6_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_7_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_7_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_7_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_7_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_7_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_7_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_7_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_7_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_7_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_7_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_7_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_8_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_8_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_8_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_8_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_8_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_8_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_8_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_8_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_8_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_8_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_8_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_9_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_9_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_9_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_9_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_9_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_9_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_9_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_9_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_9_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_9_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_9_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_10_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_10_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_10_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_10_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_10_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_10_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_10_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_10_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_10_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_10_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_10_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_11_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_11_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_11_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_11_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_11_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_11_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_11_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_11_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_11_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_11_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_11_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_12_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_12_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_12_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_12_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_12_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_12_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_12_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_12_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_12_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_12_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_12_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_13_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_13_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_13_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_13_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_13_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_13_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_13_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_13_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_13_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_13_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_13_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_14_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_14_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_14_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_14_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_14_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_14_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_14_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_14_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_14_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_14_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_14_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_15_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_15_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_15_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_15_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_15_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_15_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_15_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_15_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_15_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_15_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_15_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_16_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_16_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_16_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_16_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_16_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_16_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_16_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_16_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_16_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_16_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_16_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_17_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_17_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_17_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_17_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_17_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_17_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_17_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_17_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_17_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_17_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_17_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_18_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_18_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_18_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_18_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_18_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_18_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_18_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_18_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_18_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_18_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_18_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_19_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_19_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_19_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_19_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_19_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_19_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_19_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_19_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_19_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_19_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_19_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_20_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_20_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_20_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_20_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_20_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_20_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_20_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_20_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_20_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_20_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_20_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_21_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_21_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_21_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_21_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_21_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_21_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_21_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_21_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_21_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_21_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_21_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_22_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_22_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_22_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_22_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_22_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_22_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_22_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_22_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_22_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_22_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_22_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_23_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_23_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_23_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_23_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_23_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_23_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_23_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_23_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_23_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_23_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_23_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_24_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_24_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_24_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_24_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_24_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_24_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_24_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_24_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_24_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_24_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_24_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_25_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_25_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_25_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_25_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_25_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_25_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_25_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_25_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_25_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_25_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_25_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_26_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_26_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_26_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_26_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_26_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_26_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_26_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_26_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_26_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_26_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_26_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_27_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_27_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_27_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_27_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_27_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_27_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_27_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_27_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_27_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_27_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_27_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_28_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_28_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_28_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_28_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_28_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_28_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_28_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_28_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_28_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_28_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_28_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_29_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_29_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_29_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_29_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_29_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_29_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_29_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_29_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_29_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_29_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_29_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_30_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_30_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_30_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_30_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_30_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_30_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_30_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_30_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_30_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_30_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_30_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_31_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_31_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_31_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_31_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_31_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_31_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_31_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_31_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_31_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_31_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_31_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_32_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_32_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_32_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_32_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_32_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_32_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_32_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_32_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_32_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_32_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_32_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_33_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_33_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_33_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_33_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_33_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_33_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_33_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_33_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_33_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_33_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_33_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_34_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_34_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_34_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_34_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_34_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_34_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_34_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_34_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_34_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_34_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_34_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_35_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_35_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_35_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_35_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_35_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_35_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_35_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_35_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_35_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_35_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_35_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_36_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_36_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_36_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_36_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_36_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_36_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_36_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_36_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_36_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_36_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_36_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_37_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_37_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_37_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_37_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_37_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_37_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_37_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_37_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_37_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_37_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_37_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_38_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_38_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_38_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_38_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_38_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_38_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_38_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_38_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_38_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_38_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_38_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_39_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_39_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_39_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_39_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_39_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_39_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_39_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_39_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_39_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_39_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_39_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_40_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_40_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_40_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_40_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_40_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_40_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_40_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_40_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_40_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_40_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_40_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_41_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_41_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_41_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_41_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_41_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_41_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_41_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_41_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_41_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_41_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_41_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_42_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_42_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_42_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_42_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_42_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_42_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_42_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_42_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_42_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_42_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_42_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_43_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_43_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_43_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_43_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_43_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_43_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_43_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_43_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_43_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_43_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_43_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_44_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_44_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_44_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_44_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_44_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_44_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_44_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_44_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_44_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_44_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_44_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_45_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_45_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_45_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_45_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_45_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_45_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_45_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_45_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_45_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_45_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_45_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_46_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_46_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_46_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_46_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_46_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_46_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_46_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_46_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_46_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_46_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_46_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_47_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_47_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_47_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_47_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_47_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_47_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_47_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_47_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_47_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_47_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_47_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_48_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_48_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_48_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_48_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_48_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_48_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_48_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_48_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_48_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_48_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_48_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_49_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_49_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_49_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_49_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_49_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_49_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_49_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_49_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_49_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_49_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_49_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_50_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_50_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_50_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_50_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_50_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_50_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_50_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_50_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_50_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_50_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_50_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_51_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_51_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_51_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_51_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_51_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_51_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_51_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_51_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_51_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_51_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_51_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_52_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_52_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_52_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_52_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_52_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_52_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_52_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_52_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_52_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_52_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_52_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_53_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_53_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_53_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_53_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_53_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_53_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_53_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_53_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_53_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_53_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_53_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_54_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_54_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_54_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_54_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_54_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_54_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_54_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_54_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_54_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_54_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_54_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_55_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_55_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_55_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_55_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_55_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_55_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_55_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_55_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_55_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_55_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_55_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_56_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_56_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_56_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_56_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_56_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_56_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_56_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_56_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_56_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_56_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_56_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_57_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_57_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_57_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_57_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_57_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_57_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_57_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_57_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_57_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_57_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_57_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_58_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_58_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_58_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_58_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_58_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_58_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_58_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_58_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_58_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_58_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_58_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_59_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_59_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_59_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_59_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_59_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_59_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_59_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_59_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_59_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_59_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_59_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_60_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_60_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_60_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_60_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_60_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_60_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_60_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_60_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_60_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_60_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_60_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_61_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_61_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_61_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_61_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_61_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_61_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_61_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_61_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_61_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_61_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_61_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_62_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_62_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_62_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_62_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_62_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_62_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_62_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_62_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_62_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_62_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_62_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_63_clock; // @[contNetwork.scala 16:53]
  wire  networkUnits_63_reset; // @[contNetwork.scala 16:53]
  wire  networkUnits_63_io_addressIn_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_63_io_addressIn_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_63_io_addressIn_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_63_io_addressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_63_io_addressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_63_io_addressOut_bits; // @[contNetwork.scala 16:53]
  wire  networkUnits_63_io_casAddressOut_ready; // @[contNetwork.scala 16:53]
  wire  networkUnits_63_io_casAddressOut_valid; // @[contNetwork.scala 16:53]
  wire [63:0] networkUnits_63_io_casAddressOut_bits; // @[contNetwork.scala 16:53]
  wire  casServers_0_clock; // @[contNetwork.scala 17:53]
  wire  casServers_0_reset; // @[contNetwork.scala 17:53]
  wire  casServers_0_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_0_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_0_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_0_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_0_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_0_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_1_clock; // @[contNetwork.scala 17:53]
  wire  casServers_1_reset; // @[contNetwork.scala 17:53]
  wire  casServers_1_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_1_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_1_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_1_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_1_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_1_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_2_clock; // @[contNetwork.scala 17:53]
  wire  casServers_2_reset; // @[contNetwork.scala 17:53]
  wire  casServers_2_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_2_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_2_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_2_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_2_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_2_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_3_clock; // @[contNetwork.scala 17:53]
  wire  casServers_3_reset; // @[contNetwork.scala 17:53]
  wire  casServers_3_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_3_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_3_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_3_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_3_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_3_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_4_clock; // @[contNetwork.scala 17:53]
  wire  casServers_4_reset; // @[contNetwork.scala 17:53]
  wire  casServers_4_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_4_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_4_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_4_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_4_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_4_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_5_clock; // @[contNetwork.scala 17:53]
  wire  casServers_5_reset; // @[contNetwork.scala 17:53]
  wire  casServers_5_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_5_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_5_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_5_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_5_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_5_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_6_clock; // @[contNetwork.scala 17:53]
  wire  casServers_6_reset; // @[contNetwork.scala 17:53]
  wire  casServers_6_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_6_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_6_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_6_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_6_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_6_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_7_clock; // @[contNetwork.scala 17:53]
  wire  casServers_7_reset; // @[contNetwork.scala 17:53]
  wire  casServers_7_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_7_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_7_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_7_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_7_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_7_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_8_clock; // @[contNetwork.scala 17:53]
  wire  casServers_8_reset; // @[contNetwork.scala 17:53]
  wire  casServers_8_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_8_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_8_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_8_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_8_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_8_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_9_clock; // @[contNetwork.scala 17:53]
  wire  casServers_9_reset; // @[contNetwork.scala 17:53]
  wire  casServers_9_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_9_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_9_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_9_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_9_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_9_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_10_clock; // @[contNetwork.scala 17:53]
  wire  casServers_10_reset; // @[contNetwork.scala 17:53]
  wire  casServers_10_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_10_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_10_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_10_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_10_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_10_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_11_clock; // @[contNetwork.scala 17:53]
  wire  casServers_11_reset; // @[contNetwork.scala 17:53]
  wire  casServers_11_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_11_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_11_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_11_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_11_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_11_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_12_clock; // @[contNetwork.scala 17:53]
  wire  casServers_12_reset; // @[contNetwork.scala 17:53]
  wire  casServers_12_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_12_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_12_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_12_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_12_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_12_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_13_clock; // @[contNetwork.scala 17:53]
  wire  casServers_13_reset; // @[contNetwork.scala 17:53]
  wire  casServers_13_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_13_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_13_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_13_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_13_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_13_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_14_clock; // @[contNetwork.scala 17:53]
  wire  casServers_14_reset; // @[contNetwork.scala 17:53]
  wire  casServers_14_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_14_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_14_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_14_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_14_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_14_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_15_clock; // @[contNetwork.scala 17:53]
  wire  casServers_15_reset; // @[contNetwork.scala 17:53]
  wire  casServers_15_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_15_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_15_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_15_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_15_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_15_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_16_clock; // @[contNetwork.scala 17:53]
  wire  casServers_16_reset; // @[contNetwork.scala 17:53]
  wire  casServers_16_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_16_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_16_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_16_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_16_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_16_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_17_clock; // @[contNetwork.scala 17:53]
  wire  casServers_17_reset; // @[contNetwork.scala 17:53]
  wire  casServers_17_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_17_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_17_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_17_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_17_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_17_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_18_clock; // @[contNetwork.scala 17:53]
  wire  casServers_18_reset; // @[contNetwork.scala 17:53]
  wire  casServers_18_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_18_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_18_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_18_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_18_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_18_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_19_clock; // @[contNetwork.scala 17:53]
  wire  casServers_19_reset; // @[contNetwork.scala 17:53]
  wire  casServers_19_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_19_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_19_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_19_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_19_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_19_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_20_clock; // @[contNetwork.scala 17:53]
  wire  casServers_20_reset; // @[contNetwork.scala 17:53]
  wire  casServers_20_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_20_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_20_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_20_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_20_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_20_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_21_clock; // @[contNetwork.scala 17:53]
  wire  casServers_21_reset; // @[contNetwork.scala 17:53]
  wire  casServers_21_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_21_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_21_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_21_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_21_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_21_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_22_clock; // @[contNetwork.scala 17:53]
  wire  casServers_22_reset; // @[contNetwork.scala 17:53]
  wire  casServers_22_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_22_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_22_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_22_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_22_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_22_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_23_clock; // @[contNetwork.scala 17:53]
  wire  casServers_23_reset; // @[contNetwork.scala 17:53]
  wire  casServers_23_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_23_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_23_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_23_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_23_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_23_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_24_clock; // @[contNetwork.scala 17:53]
  wire  casServers_24_reset; // @[contNetwork.scala 17:53]
  wire  casServers_24_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_24_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_24_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_24_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_24_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_24_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_25_clock; // @[contNetwork.scala 17:53]
  wire  casServers_25_reset; // @[contNetwork.scala 17:53]
  wire  casServers_25_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_25_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_25_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_25_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_25_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_25_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_26_clock; // @[contNetwork.scala 17:53]
  wire  casServers_26_reset; // @[contNetwork.scala 17:53]
  wire  casServers_26_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_26_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_26_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_26_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_26_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_26_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_27_clock; // @[contNetwork.scala 17:53]
  wire  casServers_27_reset; // @[contNetwork.scala 17:53]
  wire  casServers_27_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_27_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_27_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_27_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_27_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_27_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_28_clock; // @[contNetwork.scala 17:53]
  wire  casServers_28_reset; // @[contNetwork.scala 17:53]
  wire  casServers_28_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_28_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_28_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_28_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_28_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_28_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_29_clock; // @[contNetwork.scala 17:53]
  wire  casServers_29_reset; // @[contNetwork.scala 17:53]
  wire  casServers_29_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_29_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_29_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_29_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_29_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_29_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_30_clock; // @[contNetwork.scala 17:53]
  wire  casServers_30_reset; // @[contNetwork.scala 17:53]
  wire  casServers_30_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_30_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_30_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_30_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_30_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_30_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_31_clock; // @[contNetwork.scala 17:53]
  wire  casServers_31_reset; // @[contNetwork.scala 17:53]
  wire  casServers_31_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_31_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_31_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_31_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_31_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_31_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_32_clock; // @[contNetwork.scala 17:53]
  wire  casServers_32_reset; // @[contNetwork.scala 17:53]
  wire  casServers_32_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_32_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_32_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_32_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_32_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_32_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_33_clock; // @[contNetwork.scala 17:53]
  wire  casServers_33_reset; // @[contNetwork.scala 17:53]
  wire  casServers_33_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_33_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_33_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_33_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_33_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_33_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_34_clock; // @[contNetwork.scala 17:53]
  wire  casServers_34_reset; // @[contNetwork.scala 17:53]
  wire  casServers_34_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_34_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_34_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_34_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_34_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_34_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_35_clock; // @[contNetwork.scala 17:53]
  wire  casServers_35_reset; // @[contNetwork.scala 17:53]
  wire  casServers_35_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_35_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_35_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_35_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_35_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_35_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_36_clock; // @[contNetwork.scala 17:53]
  wire  casServers_36_reset; // @[contNetwork.scala 17:53]
  wire  casServers_36_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_36_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_36_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_36_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_36_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_36_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_37_clock; // @[contNetwork.scala 17:53]
  wire  casServers_37_reset; // @[contNetwork.scala 17:53]
  wire  casServers_37_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_37_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_37_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_37_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_37_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_37_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_38_clock; // @[contNetwork.scala 17:53]
  wire  casServers_38_reset; // @[contNetwork.scala 17:53]
  wire  casServers_38_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_38_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_38_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_38_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_38_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_38_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_39_clock; // @[contNetwork.scala 17:53]
  wire  casServers_39_reset; // @[contNetwork.scala 17:53]
  wire  casServers_39_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_39_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_39_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_39_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_39_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_39_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_40_clock; // @[contNetwork.scala 17:53]
  wire  casServers_40_reset; // @[contNetwork.scala 17:53]
  wire  casServers_40_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_40_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_40_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_40_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_40_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_40_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_41_clock; // @[contNetwork.scala 17:53]
  wire  casServers_41_reset; // @[contNetwork.scala 17:53]
  wire  casServers_41_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_41_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_41_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_41_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_41_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_41_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_42_clock; // @[contNetwork.scala 17:53]
  wire  casServers_42_reset; // @[contNetwork.scala 17:53]
  wire  casServers_42_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_42_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_42_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_42_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_42_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_42_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_43_clock; // @[contNetwork.scala 17:53]
  wire  casServers_43_reset; // @[contNetwork.scala 17:53]
  wire  casServers_43_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_43_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_43_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_43_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_43_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_43_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_44_clock; // @[contNetwork.scala 17:53]
  wire  casServers_44_reset; // @[contNetwork.scala 17:53]
  wire  casServers_44_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_44_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_44_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_44_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_44_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_44_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_45_clock; // @[contNetwork.scala 17:53]
  wire  casServers_45_reset; // @[contNetwork.scala 17:53]
  wire  casServers_45_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_45_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_45_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_45_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_45_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_45_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_46_clock; // @[contNetwork.scala 17:53]
  wire  casServers_46_reset; // @[contNetwork.scala 17:53]
  wire  casServers_46_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_46_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_46_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_46_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_46_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_46_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_47_clock; // @[contNetwork.scala 17:53]
  wire  casServers_47_reset; // @[contNetwork.scala 17:53]
  wire  casServers_47_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_47_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_47_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_47_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_47_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_47_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_48_clock; // @[contNetwork.scala 17:53]
  wire  casServers_48_reset; // @[contNetwork.scala 17:53]
  wire  casServers_48_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_48_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_48_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_48_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_48_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_48_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_49_clock; // @[contNetwork.scala 17:53]
  wire  casServers_49_reset; // @[contNetwork.scala 17:53]
  wire  casServers_49_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_49_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_49_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_49_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_49_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_49_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_50_clock; // @[contNetwork.scala 17:53]
  wire  casServers_50_reset; // @[contNetwork.scala 17:53]
  wire  casServers_50_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_50_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_50_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_50_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_50_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_50_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_51_clock; // @[contNetwork.scala 17:53]
  wire  casServers_51_reset; // @[contNetwork.scala 17:53]
  wire  casServers_51_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_51_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_51_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_51_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_51_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_51_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_52_clock; // @[contNetwork.scala 17:53]
  wire  casServers_52_reset; // @[contNetwork.scala 17:53]
  wire  casServers_52_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_52_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_52_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_52_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_52_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_52_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_53_clock; // @[contNetwork.scala 17:53]
  wire  casServers_53_reset; // @[contNetwork.scala 17:53]
  wire  casServers_53_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_53_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_53_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_53_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_53_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_53_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_54_clock; // @[contNetwork.scala 17:53]
  wire  casServers_54_reset; // @[contNetwork.scala 17:53]
  wire  casServers_54_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_54_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_54_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_54_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_54_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_54_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_55_clock; // @[contNetwork.scala 17:53]
  wire  casServers_55_reset; // @[contNetwork.scala 17:53]
  wire  casServers_55_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_55_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_55_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_55_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_55_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_55_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_56_clock; // @[contNetwork.scala 17:53]
  wire  casServers_56_reset; // @[contNetwork.scala 17:53]
  wire  casServers_56_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_56_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_56_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_56_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_56_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_56_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_57_clock; // @[contNetwork.scala 17:53]
  wire  casServers_57_reset; // @[contNetwork.scala 17:53]
  wire  casServers_57_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_57_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_57_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_57_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_57_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_57_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_58_clock; // @[contNetwork.scala 17:53]
  wire  casServers_58_reset; // @[contNetwork.scala 17:53]
  wire  casServers_58_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_58_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_58_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_58_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_58_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_58_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_59_clock; // @[contNetwork.scala 17:53]
  wire  casServers_59_reset; // @[contNetwork.scala 17:53]
  wire  casServers_59_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_59_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_59_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_59_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_59_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_59_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_60_clock; // @[contNetwork.scala 17:53]
  wire  casServers_60_reset; // @[contNetwork.scala 17:53]
  wire  casServers_60_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_60_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_60_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_60_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_60_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_60_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_61_clock; // @[contNetwork.scala 17:53]
  wire  casServers_61_reset; // @[contNetwork.scala 17:53]
  wire  casServers_61_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_61_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_61_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_61_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_61_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_61_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_62_clock; // @[contNetwork.scala 17:53]
  wire  casServers_62_reset; // @[contNetwork.scala 17:53]
  wire  casServers_62_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_62_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_62_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_62_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_62_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_62_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  casServers_63_clock; // @[contNetwork.scala 17:53]
  wire  casServers_63_reset; // @[contNetwork.scala 17:53]
  wire  casServers_63_io_addressIn_ready; // @[contNetwork.scala 17:53]
  wire  casServers_63_io_addressIn_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_63_io_addressIn_bits; // @[contNetwork.scala 17:53]
  wire  casServers_63_io_addressOut_ready; // @[contNetwork.scala 17:53]
  wire  casServers_63_io_addressOut_valid; // @[contNetwork.scala 17:53]
  wire [63:0] casServers_63_io_addressOut_bits; // @[contNetwork.scala 17:53]
  wire  queues_0_clock; // @[contNetwork.scala 18:53]
  wire  queues_0_reset; // @[contNetwork.scala 18:53]
  wire  queues_0_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_0_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_0_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_0_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_0_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_0_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_1_clock; // @[contNetwork.scala 18:53]
  wire  queues_1_reset; // @[contNetwork.scala 18:53]
  wire  queues_1_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_1_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_1_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_1_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_1_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_1_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_2_clock; // @[contNetwork.scala 18:53]
  wire  queues_2_reset; // @[contNetwork.scala 18:53]
  wire  queues_2_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_2_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_2_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_2_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_2_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_2_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_3_clock; // @[contNetwork.scala 18:53]
  wire  queues_3_reset; // @[contNetwork.scala 18:53]
  wire  queues_3_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_3_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_3_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_3_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_3_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_3_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_4_clock; // @[contNetwork.scala 18:53]
  wire  queues_4_reset; // @[contNetwork.scala 18:53]
  wire  queues_4_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_4_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_4_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_4_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_4_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_4_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_5_clock; // @[contNetwork.scala 18:53]
  wire  queues_5_reset; // @[contNetwork.scala 18:53]
  wire  queues_5_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_5_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_5_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_5_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_5_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_5_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_6_clock; // @[contNetwork.scala 18:53]
  wire  queues_6_reset; // @[contNetwork.scala 18:53]
  wire  queues_6_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_6_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_6_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_6_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_6_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_6_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_7_clock; // @[contNetwork.scala 18:53]
  wire  queues_7_reset; // @[contNetwork.scala 18:53]
  wire  queues_7_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_7_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_7_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_7_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_7_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_7_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_8_clock; // @[contNetwork.scala 18:53]
  wire  queues_8_reset; // @[contNetwork.scala 18:53]
  wire  queues_8_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_8_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_8_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_8_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_8_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_8_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_9_clock; // @[contNetwork.scala 18:53]
  wire  queues_9_reset; // @[contNetwork.scala 18:53]
  wire  queues_9_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_9_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_9_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_9_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_9_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_9_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_10_clock; // @[contNetwork.scala 18:53]
  wire  queues_10_reset; // @[contNetwork.scala 18:53]
  wire  queues_10_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_10_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_10_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_10_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_10_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_10_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_11_clock; // @[contNetwork.scala 18:53]
  wire  queues_11_reset; // @[contNetwork.scala 18:53]
  wire  queues_11_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_11_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_11_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_11_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_11_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_11_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_12_clock; // @[contNetwork.scala 18:53]
  wire  queues_12_reset; // @[contNetwork.scala 18:53]
  wire  queues_12_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_12_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_12_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_12_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_12_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_12_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_13_clock; // @[contNetwork.scala 18:53]
  wire  queues_13_reset; // @[contNetwork.scala 18:53]
  wire  queues_13_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_13_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_13_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_13_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_13_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_13_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_14_clock; // @[contNetwork.scala 18:53]
  wire  queues_14_reset; // @[contNetwork.scala 18:53]
  wire  queues_14_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_14_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_14_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_14_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_14_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_14_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_15_clock; // @[contNetwork.scala 18:53]
  wire  queues_15_reset; // @[contNetwork.scala 18:53]
  wire  queues_15_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_15_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_15_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_15_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_15_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_15_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_16_clock; // @[contNetwork.scala 18:53]
  wire  queues_16_reset; // @[contNetwork.scala 18:53]
  wire  queues_16_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_16_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_16_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_16_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_16_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_16_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_17_clock; // @[contNetwork.scala 18:53]
  wire  queues_17_reset; // @[contNetwork.scala 18:53]
  wire  queues_17_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_17_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_17_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_17_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_17_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_17_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_18_clock; // @[contNetwork.scala 18:53]
  wire  queues_18_reset; // @[contNetwork.scala 18:53]
  wire  queues_18_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_18_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_18_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_18_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_18_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_18_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_19_clock; // @[contNetwork.scala 18:53]
  wire  queues_19_reset; // @[contNetwork.scala 18:53]
  wire  queues_19_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_19_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_19_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_19_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_19_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_19_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_20_clock; // @[contNetwork.scala 18:53]
  wire  queues_20_reset; // @[contNetwork.scala 18:53]
  wire  queues_20_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_20_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_20_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_20_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_20_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_20_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_21_clock; // @[contNetwork.scala 18:53]
  wire  queues_21_reset; // @[contNetwork.scala 18:53]
  wire  queues_21_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_21_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_21_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_21_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_21_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_21_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_22_clock; // @[contNetwork.scala 18:53]
  wire  queues_22_reset; // @[contNetwork.scala 18:53]
  wire  queues_22_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_22_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_22_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_22_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_22_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_22_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_23_clock; // @[contNetwork.scala 18:53]
  wire  queues_23_reset; // @[contNetwork.scala 18:53]
  wire  queues_23_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_23_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_23_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_23_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_23_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_23_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_24_clock; // @[contNetwork.scala 18:53]
  wire  queues_24_reset; // @[contNetwork.scala 18:53]
  wire  queues_24_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_24_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_24_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_24_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_24_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_24_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_25_clock; // @[contNetwork.scala 18:53]
  wire  queues_25_reset; // @[contNetwork.scala 18:53]
  wire  queues_25_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_25_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_25_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_25_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_25_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_25_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_26_clock; // @[contNetwork.scala 18:53]
  wire  queues_26_reset; // @[contNetwork.scala 18:53]
  wire  queues_26_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_26_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_26_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_26_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_26_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_26_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_27_clock; // @[contNetwork.scala 18:53]
  wire  queues_27_reset; // @[contNetwork.scala 18:53]
  wire  queues_27_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_27_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_27_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_27_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_27_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_27_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_28_clock; // @[contNetwork.scala 18:53]
  wire  queues_28_reset; // @[contNetwork.scala 18:53]
  wire  queues_28_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_28_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_28_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_28_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_28_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_28_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_29_clock; // @[contNetwork.scala 18:53]
  wire  queues_29_reset; // @[contNetwork.scala 18:53]
  wire  queues_29_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_29_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_29_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_29_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_29_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_29_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_30_clock; // @[contNetwork.scala 18:53]
  wire  queues_30_reset; // @[contNetwork.scala 18:53]
  wire  queues_30_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_30_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_30_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_30_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_30_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_30_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_31_clock; // @[contNetwork.scala 18:53]
  wire  queues_31_reset; // @[contNetwork.scala 18:53]
  wire  queues_31_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_31_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_31_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_31_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_31_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_31_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_32_clock; // @[contNetwork.scala 18:53]
  wire  queues_32_reset; // @[contNetwork.scala 18:53]
  wire  queues_32_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_32_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_32_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_32_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_32_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_32_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_33_clock; // @[contNetwork.scala 18:53]
  wire  queues_33_reset; // @[contNetwork.scala 18:53]
  wire  queues_33_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_33_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_33_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_33_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_33_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_33_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_34_clock; // @[contNetwork.scala 18:53]
  wire  queues_34_reset; // @[contNetwork.scala 18:53]
  wire  queues_34_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_34_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_34_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_34_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_34_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_34_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_35_clock; // @[contNetwork.scala 18:53]
  wire  queues_35_reset; // @[contNetwork.scala 18:53]
  wire  queues_35_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_35_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_35_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_35_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_35_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_35_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_36_clock; // @[contNetwork.scala 18:53]
  wire  queues_36_reset; // @[contNetwork.scala 18:53]
  wire  queues_36_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_36_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_36_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_36_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_36_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_36_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_37_clock; // @[contNetwork.scala 18:53]
  wire  queues_37_reset; // @[contNetwork.scala 18:53]
  wire  queues_37_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_37_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_37_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_37_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_37_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_37_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_38_clock; // @[contNetwork.scala 18:53]
  wire  queues_38_reset; // @[contNetwork.scala 18:53]
  wire  queues_38_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_38_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_38_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_38_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_38_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_38_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_39_clock; // @[contNetwork.scala 18:53]
  wire  queues_39_reset; // @[contNetwork.scala 18:53]
  wire  queues_39_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_39_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_39_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_39_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_39_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_39_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_40_clock; // @[contNetwork.scala 18:53]
  wire  queues_40_reset; // @[contNetwork.scala 18:53]
  wire  queues_40_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_40_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_40_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_40_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_40_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_40_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_41_clock; // @[contNetwork.scala 18:53]
  wire  queues_41_reset; // @[contNetwork.scala 18:53]
  wire  queues_41_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_41_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_41_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_41_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_41_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_41_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_42_clock; // @[contNetwork.scala 18:53]
  wire  queues_42_reset; // @[contNetwork.scala 18:53]
  wire  queues_42_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_42_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_42_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_42_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_42_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_42_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_43_clock; // @[contNetwork.scala 18:53]
  wire  queues_43_reset; // @[contNetwork.scala 18:53]
  wire  queues_43_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_43_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_43_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_43_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_43_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_43_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_44_clock; // @[contNetwork.scala 18:53]
  wire  queues_44_reset; // @[contNetwork.scala 18:53]
  wire  queues_44_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_44_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_44_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_44_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_44_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_44_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_45_clock; // @[contNetwork.scala 18:53]
  wire  queues_45_reset; // @[contNetwork.scala 18:53]
  wire  queues_45_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_45_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_45_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_45_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_45_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_45_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_46_clock; // @[contNetwork.scala 18:53]
  wire  queues_46_reset; // @[contNetwork.scala 18:53]
  wire  queues_46_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_46_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_46_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_46_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_46_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_46_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_47_clock; // @[contNetwork.scala 18:53]
  wire  queues_47_reset; // @[contNetwork.scala 18:53]
  wire  queues_47_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_47_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_47_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_47_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_47_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_47_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_48_clock; // @[contNetwork.scala 18:53]
  wire  queues_48_reset; // @[contNetwork.scala 18:53]
  wire  queues_48_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_48_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_48_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_48_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_48_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_48_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_49_clock; // @[contNetwork.scala 18:53]
  wire  queues_49_reset; // @[contNetwork.scala 18:53]
  wire  queues_49_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_49_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_49_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_49_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_49_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_49_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_50_clock; // @[contNetwork.scala 18:53]
  wire  queues_50_reset; // @[contNetwork.scala 18:53]
  wire  queues_50_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_50_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_50_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_50_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_50_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_50_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_51_clock; // @[contNetwork.scala 18:53]
  wire  queues_51_reset; // @[contNetwork.scala 18:53]
  wire  queues_51_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_51_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_51_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_51_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_51_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_51_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_52_clock; // @[contNetwork.scala 18:53]
  wire  queues_52_reset; // @[contNetwork.scala 18:53]
  wire  queues_52_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_52_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_52_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_52_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_52_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_52_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_53_clock; // @[contNetwork.scala 18:53]
  wire  queues_53_reset; // @[contNetwork.scala 18:53]
  wire  queues_53_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_53_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_53_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_53_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_53_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_53_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_54_clock; // @[contNetwork.scala 18:53]
  wire  queues_54_reset; // @[contNetwork.scala 18:53]
  wire  queues_54_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_54_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_54_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_54_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_54_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_54_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_55_clock; // @[contNetwork.scala 18:53]
  wire  queues_55_reset; // @[contNetwork.scala 18:53]
  wire  queues_55_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_55_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_55_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_55_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_55_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_55_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_56_clock; // @[contNetwork.scala 18:53]
  wire  queues_56_reset; // @[contNetwork.scala 18:53]
  wire  queues_56_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_56_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_56_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_56_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_56_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_56_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_57_clock; // @[contNetwork.scala 18:53]
  wire  queues_57_reset; // @[contNetwork.scala 18:53]
  wire  queues_57_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_57_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_57_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_57_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_57_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_57_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_58_clock; // @[contNetwork.scala 18:53]
  wire  queues_58_reset; // @[contNetwork.scala 18:53]
  wire  queues_58_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_58_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_58_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_58_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_58_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_58_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_59_clock; // @[contNetwork.scala 18:53]
  wire  queues_59_reset; // @[contNetwork.scala 18:53]
  wire  queues_59_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_59_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_59_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_59_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_59_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_59_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_60_clock; // @[contNetwork.scala 18:53]
  wire  queues_60_reset; // @[contNetwork.scala 18:53]
  wire  queues_60_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_60_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_60_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_60_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_60_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_60_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_61_clock; // @[contNetwork.scala 18:53]
  wire  queues_61_reset; // @[contNetwork.scala 18:53]
  wire  queues_61_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_61_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_61_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_61_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_61_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_61_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_62_clock; // @[contNetwork.scala 18:53]
  wire  queues_62_reset; // @[contNetwork.scala 18:53]
  wire  queues_62_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_62_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_62_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_62_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_62_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_62_io_addressOut_bits; // @[contNetwork.scala 18:53]
  wire  queues_63_clock; // @[contNetwork.scala 18:53]
  wire  queues_63_reset; // @[contNetwork.scala 18:53]
  wire  queues_63_io_addressIn_ready; // @[contNetwork.scala 18:53]
  wire  queues_63_io_addressIn_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_63_io_addressIn_bits; // @[contNetwork.scala 18:53]
  wire  queues_63_io_addressOut_ready; // @[contNetwork.scala 18:53]
  wire  queues_63_io_addressOut_valid; // @[contNetwork.scala 18:53]
  wire [63:0] queues_63_io_addressOut_bits; // @[contNetwork.scala 18:53]
  contAddrNtwUnitCAS vcasNetworkUnits_0 ( // @[contNetwork.scala 15:55]
    .clock(vcasNetworkUnits_0_clock),
    .reset(vcasNetworkUnits_0_reset),
    .io_addressIn1_ready(vcasNetworkUnits_0_io_addressIn1_ready),
    .io_addressIn1_valid(vcasNetworkUnits_0_io_addressIn1_valid),
    .io_addressIn1_bits(vcasNetworkUnits_0_io_addressIn1_bits),
    .io_addressOut_ready(vcasNetworkUnits_0_io_addressOut_ready),
    .io_addressOut_valid(vcasNetworkUnits_0_io_addressOut_valid),
    .io_addressOut_bits(vcasNetworkUnits_0_io_addressOut_bits)
  );
  contAddrNtwUnit networkUnits_0 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_0_clock),
    .reset(networkUnits_0_reset),
    .io_addressIn_ready(networkUnits_0_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_0_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_0_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_0_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_0_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_0_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_0_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_0_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_0_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_1 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_1_clock),
    .reset(networkUnits_1_reset),
    .io_addressIn_ready(networkUnits_1_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_1_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_1_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_1_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_1_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_1_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_1_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_1_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_1_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_2 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_2_clock),
    .reset(networkUnits_2_reset),
    .io_addressIn_ready(networkUnits_2_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_2_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_2_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_2_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_2_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_2_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_2_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_2_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_2_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_3 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_3_clock),
    .reset(networkUnits_3_reset),
    .io_addressIn_ready(networkUnits_3_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_3_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_3_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_3_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_3_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_3_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_3_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_3_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_3_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_4 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_4_clock),
    .reset(networkUnits_4_reset),
    .io_addressIn_ready(networkUnits_4_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_4_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_4_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_4_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_4_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_4_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_4_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_4_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_4_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_5 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_5_clock),
    .reset(networkUnits_5_reset),
    .io_addressIn_ready(networkUnits_5_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_5_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_5_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_5_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_5_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_5_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_5_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_5_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_5_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_6 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_6_clock),
    .reset(networkUnits_6_reset),
    .io_addressIn_ready(networkUnits_6_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_6_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_6_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_6_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_6_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_6_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_6_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_6_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_6_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_7 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_7_clock),
    .reset(networkUnits_7_reset),
    .io_addressIn_ready(networkUnits_7_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_7_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_7_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_7_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_7_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_7_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_7_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_7_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_7_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_8 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_8_clock),
    .reset(networkUnits_8_reset),
    .io_addressIn_ready(networkUnits_8_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_8_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_8_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_8_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_8_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_8_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_8_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_8_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_8_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_9 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_9_clock),
    .reset(networkUnits_9_reset),
    .io_addressIn_ready(networkUnits_9_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_9_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_9_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_9_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_9_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_9_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_9_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_9_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_9_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_10 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_10_clock),
    .reset(networkUnits_10_reset),
    .io_addressIn_ready(networkUnits_10_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_10_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_10_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_10_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_10_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_10_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_10_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_10_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_10_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_11 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_11_clock),
    .reset(networkUnits_11_reset),
    .io_addressIn_ready(networkUnits_11_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_11_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_11_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_11_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_11_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_11_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_11_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_11_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_11_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_12 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_12_clock),
    .reset(networkUnits_12_reset),
    .io_addressIn_ready(networkUnits_12_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_12_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_12_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_12_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_12_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_12_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_12_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_12_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_12_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_13 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_13_clock),
    .reset(networkUnits_13_reset),
    .io_addressIn_ready(networkUnits_13_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_13_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_13_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_13_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_13_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_13_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_13_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_13_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_13_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_14 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_14_clock),
    .reset(networkUnits_14_reset),
    .io_addressIn_ready(networkUnits_14_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_14_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_14_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_14_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_14_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_14_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_14_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_14_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_14_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_15 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_15_clock),
    .reset(networkUnits_15_reset),
    .io_addressIn_ready(networkUnits_15_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_15_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_15_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_15_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_15_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_15_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_15_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_15_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_15_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_16 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_16_clock),
    .reset(networkUnits_16_reset),
    .io_addressIn_ready(networkUnits_16_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_16_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_16_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_16_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_16_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_16_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_16_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_16_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_16_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_17 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_17_clock),
    .reset(networkUnits_17_reset),
    .io_addressIn_ready(networkUnits_17_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_17_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_17_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_17_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_17_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_17_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_17_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_17_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_17_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_18 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_18_clock),
    .reset(networkUnits_18_reset),
    .io_addressIn_ready(networkUnits_18_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_18_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_18_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_18_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_18_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_18_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_18_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_18_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_18_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_19 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_19_clock),
    .reset(networkUnits_19_reset),
    .io_addressIn_ready(networkUnits_19_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_19_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_19_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_19_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_19_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_19_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_19_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_19_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_19_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_20 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_20_clock),
    .reset(networkUnits_20_reset),
    .io_addressIn_ready(networkUnits_20_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_20_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_20_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_20_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_20_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_20_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_20_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_20_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_20_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_21 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_21_clock),
    .reset(networkUnits_21_reset),
    .io_addressIn_ready(networkUnits_21_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_21_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_21_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_21_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_21_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_21_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_21_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_21_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_21_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_22 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_22_clock),
    .reset(networkUnits_22_reset),
    .io_addressIn_ready(networkUnits_22_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_22_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_22_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_22_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_22_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_22_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_22_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_22_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_22_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_23 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_23_clock),
    .reset(networkUnits_23_reset),
    .io_addressIn_ready(networkUnits_23_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_23_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_23_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_23_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_23_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_23_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_23_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_23_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_23_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_24 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_24_clock),
    .reset(networkUnits_24_reset),
    .io_addressIn_ready(networkUnits_24_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_24_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_24_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_24_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_24_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_24_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_24_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_24_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_24_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_25 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_25_clock),
    .reset(networkUnits_25_reset),
    .io_addressIn_ready(networkUnits_25_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_25_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_25_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_25_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_25_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_25_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_25_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_25_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_25_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_26 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_26_clock),
    .reset(networkUnits_26_reset),
    .io_addressIn_ready(networkUnits_26_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_26_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_26_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_26_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_26_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_26_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_26_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_26_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_26_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_27 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_27_clock),
    .reset(networkUnits_27_reset),
    .io_addressIn_ready(networkUnits_27_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_27_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_27_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_27_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_27_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_27_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_27_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_27_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_27_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_28 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_28_clock),
    .reset(networkUnits_28_reset),
    .io_addressIn_ready(networkUnits_28_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_28_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_28_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_28_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_28_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_28_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_28_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_28_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_28_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_29 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_29_clock),
    .reset(networkUnits_29_reset),
    .io_addressIn_ready(networkUnits_29_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_29_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_29_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_29_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_29_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_29_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_29_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_29_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_29_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_30 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_30_clock),
    .reset(networkUnits_30_reset),
    .io_addressIn_ready(networkUnits_30_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_30_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_30_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_30_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_30_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_30_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_30_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_30_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_30_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_31 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_31_clock),
    .reset(networkUnits_31_reset),
    .io_addressIn_ready(networkUnits_31_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_31_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_31_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_31_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_31_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_31_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_31_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_31_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_31_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_32 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_32_clock),
    .reset(networkUnits_32_reset),
    .io_addressIn_ready(networkUnits_32_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_32_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_32_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_32_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_32_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_32_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_32_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_32_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_32_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_33 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_33_clock),
    .reset(networkUnits_33_reset),
    .io_addressIn_ready(networkUnits_33_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_33_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_33_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_33_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_33_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_33_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_33_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_33_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_33_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_34 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_34_clock),
    .reset(networkUnits_34_reset),
    .io_addressIn_ready(networkUnits_34_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_34_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_34_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_34_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_34_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_34_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_34_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_34_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_34_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_35 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_35_clock),
    .reset(networkUnits_35_reset),
    .io_addressIn_ready(networkUnits_35_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_35_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_35_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_35_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_35_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_35_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_35_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_35_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_35_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_36 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_36_clock),
    .reset(networkUnits_36_reset),
    .io_addressIn_ready(networkUnits_36_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_36_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_36_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_36_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_36_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_36_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_36_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_36_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_36_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_37 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_37_clock),
    .reset(networkUnits_37_reset),
    .io_addressIn_ready(networkUnits_37_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_37_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_37_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_37_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_37_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_37_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_37_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_37_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_37_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_38 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_38_clock),
    .reset(networkUnits_38_reset),
    .io_addressIn_ready(networkUnits_38_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_38_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_38_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_38_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_38_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_38_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_38_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_38_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_38_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_39 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_39_clock),
    .reset(networkUnits_39_reset),
    .io_addressIn_ready(networkUnits_39_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_39_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_39_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_39_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_39_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_39_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_39_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_39_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_39_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_40 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_40_clock),
    .reset(networkUnits_40_reset),
    .io_addressIn_ready(networkUnits_40_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_40_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_40_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_40_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_40_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_40_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_40_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_40_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_40_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_41 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_41_clock),
    .reset(networkUnits_41_reset),
    .io_addressIn_ready(networkUnits_41_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_41_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_41_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_41_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_41_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_41_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_41_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_41_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_41_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_42 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_42_clock),
    .reset(networkUnits_42_reset),
    .io_addressIn_ready(networkUnits_42_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_42_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_42_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_42_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_42_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_42_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_42_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_42_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_42_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_43 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_43_clock),
    .reset(networkUnits_43_reset),
    .io_addressIn_ready(networkUnits_43_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_43_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_43_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_43_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_43_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_43_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_43_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_43_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_43_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_44 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_44_clock),
    .reset(networkUnits_44_reset),
    .io_addressIn_ready(networkUnits_44_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_44_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_44_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_44_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_44_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_44_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_44_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_44_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_44_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_45 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_45_clock),
    .reset(networkUnits_45_reset),
    .io_addressIn_ready(networkUnits_45_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_45_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_45_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_45_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_45_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_45_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_45_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_45_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_45_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_46 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_46_clock),
    .reset(networkUnits_46_reset),
    .io_addressIn_ready(networkUnits_46_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_46_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_46_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_46_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_46_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_46_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_46_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_46_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_46_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_47 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_47_clock),
    .reset(networkUnits_47_reset),
    .io_addressIn_ready(networkUnits_47_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_47_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_47_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_47_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_47_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_47_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_47_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_47_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_47_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_48 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_48_clock),
    .reset(networkUnits_48_reset),
    .io_addressIn_ready(networkUnits_48_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_48_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_48_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_48_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_48_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_48_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_48_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_48_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_48_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_49 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_49_clock),
    .reset(networkUnits_49_reset),
    .io_addressIn_ready(networkUnits_49_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_49_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_49_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_49_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_49_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_49_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_49_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_49_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_49_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_50 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_50_clock),
    .reset(networkUnits_50_reset),
    .io_addressIn_ready(networkUnits_50_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_50_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_50_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_50_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_50_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_50_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_50_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_50_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_50_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_51 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_51_clock),
    .reset(networkUnits_51_reset),
    .io_addressIn_ready(networkUnits_51_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_51_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_51_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_51_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_51_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_51_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_51_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_51_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_51_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_52 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_52_clock),
    .reset(networkUnits_52_reset),
    .io_addressIn_ready(networkUnits_52_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_52_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_52_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_52_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_52_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_52_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_52_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_52_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_52_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_53 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_53_clock),
    .reset(networkUnits_53_reset),
    .io_addressIn_ready(networkUnits_53_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_53_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_53_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_53_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_53_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_53_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_53_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_53_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_53_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_54 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_54_clock),
    .reset(networkUnits_54_reset),
    .io_addressIn_ready(networkUnits_54_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_54_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_54_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_54_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_54_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_54_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_54_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_54_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_54_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_55 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_55_clock),
    .reset(networkUnits_55_reset),
    .io_addressIn_ready(networkUnits_55_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_55_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_55_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_55_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_55_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_55_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_55_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_55_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_55_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_56 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_56_clock),
    .reset(networkUnits_56_reset),
    .io_addressIn_ready(networkUnits_56_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_56_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_56_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_56_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_56_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_56_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_56_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_56_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_56_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_57 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_57_clock),
    .reset(networkUnits_57_reset),
    .io_addressIn_ready(networkUnits_57_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_57_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_57_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_57_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_57_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_57_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_57_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_57_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_57_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_58 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_58_clock),
    .reset(networkUnits_58_reset),
    .io_addressIn_ready(networkUnits_58_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_58_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_58_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_58_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_58_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_58_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_58_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_58_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_58_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_59 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_59_clock),
    .reset(networkUnits_59_reset),
    .io_addressIn_ready(networkUnits_59_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_59_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_59_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_59_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_59_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_59_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_59_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_59_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_59_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_60 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_60_clock),
    .reset(networkUnits_60_reset),
    .io_addressIn_ready(networkUnits_60_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_60_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_60_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_60_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_60_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_60_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_60_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_60_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_60_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_61 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_61_clock),
    .reset(networkUnits_61_reset),
    .io_addressIn_ready(networkUnits_61_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_61_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_61_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_61_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_61_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_61_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_61_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_61_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_61_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_62 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_62_clock),
    .reset(networkUnits_62_reset),
    .io_addressIn_ready(networkUnits_62_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_62_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_62_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_62_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_62_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_62_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_62_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_62_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_62_io_casAddressOut_bits)
  );
  contAddrNtwUnit networkUnits_63 ( // @[contNetwork.scala 16:53]
    .clock(networkUnits_63_clock),
    .reset(networkUnits_63_reset),
    .io_addressIn_ready(networkUnits_63_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_63_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_63_io_addressIn_bits),
    .io_addressOut_ready(networkUnits_63_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_63_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_63_io_addressOut_bits),
    .io_casAddressOut_ready(networkUnits_63_io_casAddressOut_ready),
    .io_casAddressOut_valid(networkUnits_63_io_casAddressOut_valid),
    .io_casAddressOut_bits(networkUnits_63_io_casAddressOut_bits)
  );
  contAddrServer casServers_0 ( // @[contNetwork.scala 17:53]
    .clock(casServers_0_clock),
    .reset(casServers_0_reset),
    .io_addressIn_ready(casServers_0_io_addressIn_ready),
    .io_addressIn_valid(casServers_0_io_addressIn_valid),
    .io_addressIn_bits(casServers_0_io_addressIn_bits),
    .io_addressOut_ready(casServers_0_io_addressOut_ready),
    .io_addressOut_valid(casServers_0_io_addressOut_valid),
    .io_addressOut_bits(casServers_0_io_addressOut_bits)
  );
  contAddrServer casServers_1 ( // @[contNetwork.scala 17:53]
    .clock(casServers_1_clock),
    .reset(casServers_1_reset),
    .io_addressIn_ready(casServers_1_io_addressIn_ready),
    .io_addressIn_valid(casServers_1_io_addressIn_valid),
    .io_addressIn_bits(casServers_1_io_addressIn_bits),
    .io_addressOut_ready(casServers_1_io_addressOut_ready),
    .io_addressOut_valid(casServers_1_io_addressOut_valid),
    .io_addressOut_bits(casServers_1_io_addressOut_bits)
  );
  contAddrServer casServers_2 ( // @[contNetwork.scala 17:53]
    .clock(casServers_2_clock),
    .reset(casServers_2_reset),
    .io_addressIn_ready(casServers_2_io_addressIn_ready),
    .io_addressIn_valid(casServers_2_io_addressIn_valid),
    .io_addressIn_bits(casServers_2_io_addressIn_bits),
    .io_addressOut_ready(casServers_2_io_addressOut_ready),
    .io_addressOut_valid(casServers_2_io_addressOut_valid),
    .io_addressOut_bits(casServers_2_io_addressOut_bits)
  );
  contAddrServer casServers_3 ( // @[contNetwork.scala 17:53]
    .clock(casServers_3_clock),
    .reset(casServers_3_reset),
    .io_addressIn_ready(casServers_3_io_addressIn_ready),
    .io_addressIn_valid(casServers_3_io_addressIn_valid),
    .io_addressIn_bits(casServers_3_io_addressIn_bits),
    .io_addressOut_ready(casServers_3_io_addressOut_ready),
    .io_addressOut_valid(casServers_3_io_addressOut_valid),
    .io_addressOut_bits(casServers_3_io_addressOut_bits)
  );
  contAddrServer casServers_4 ( // @[contNetwork.scala 17:53]
    .clock(casServers_4_clock),
    .reset(casServers_4_reset),
    .io_addressIn_ready(casServers_4_io_addressIn_ready),
    .io_addressIn_valid(casServers_4_io_addressIn_valid),
    .io_addressIn_bits(casServers_4_io_addressIn_bits),
    .io_addressOut_ready(casServers_4_io_addressOut_ready),
    .io_addressOut_valid(casServers_4_io_addressOut_valid),
    .io_addressOut_bits(casServers_4_io_addressOut_bits)
  );
  contAddrServer casServers_5 ( // @[contNetwork.scala 17:53]
    .clock(casServers_5_clock),
    .reset(casServers_5_reset),
    .io_addressIn_ready(casServers_5_io_addressIn_ready),
    .io_addressIn_valid(casServers_5_io_addressIn_valid),
    .io_addressIn_bits(casServers_5_io_addressIn_bits),
    .io_addressOut_ready(casServers_5_io_addressOut_ready),
    .io_addressOut_valid(casServers_5_io_addressOut_valid),
    .io_addressOut_bits(casServers_5_io_addressOut_bits)
  );
  contAddrServer casServers_6 ( // @[contNetwork.scala 17:53]
    .clock(casServers_6_clock),
    .reset(casServers_6_reset),
    .io_addressIn_ready(casServers_6_io_addressIn_ready),
    .io_addressIn_valid(casServers_6_io_addressIn_valid),
    .io_addressIn_bits(casServers_6_io_addressIn_bits),
    .io_addressOut_ready(casServers_6_io_addressOut_ready),
    .io_addressOut_valid(casServers_6_io_addressOut_valid),
    .io_addressOut_bits(casServers_6_io_addressOut_bits)
  );
  contAddrServer casServers_7 ( // @[contNetwork.scala 17:53]
    .clock(casServers_7_clock),
    .reset(casServers_7_reset),
    .io_addressIn_ready(casServers_7_io_addressIn_ready),
    .io_addressIn_valid(casServers_7_io_addressIn_valid),
    .io_addressIn_bits(casServers_7_io_addressIn_bits),
    .io_addressOut_ready(casServers_7_io_addressOut_ready),
    .io_addressOut_valid(casServers_7_io_addressOut_valid),
    .io_addressOut_bits(casServers_7_io_addressOut_bits)
  );
  contAddrServer casServers_8 ( // @[contNetwork.scala 17:53]
    .clock(casServers_8_clock),
    .reset(casServers_8_reset),
    .io_addressIn_ready(casServers_8_io_addressIn_ready),
    .io_addressIn_valid(casServers_8_io_addressIn_valid),
    .io_addressIn_bits(casServers_8_io_addressIn_bits),
    .io_addressOut_ready(casServers_8_io_addressOut_ready),
    .io_addressOut_valid(casServers_8_io_addressOut_valid),
    .io_addressOut_bits(casServers_8_io_addressOut_bits)
  );
  contAddrServer casServers_9 ( // @[contNetwork.scala 17:53]
    .clock(casServers_9_clock),
    .reset(casServers_9_reset),
    .io_addressIn_ready(casServers_9_io_addressIn_ready),
    .io_addressIn_valid(casServers_9_io_addressIn_valid),
    .io_addressIn_bits(casServers_9_io_addressIn_bits),
    .io_addressOut_ready(casServers_9_io_addressOut_ready),
    .io_addressOut_valid(casServers_9_io_addressOut_valid),
    .io_addressOut_bits(casServers_9_io_addressOut_bits)
  );
  contAddrServer casServers_10 ( // @[contNetwork.scala 17:53]
    .clock(casServers_10_clock),
    .reset(casServers_10_reset),
    .io_addressIn_ready(casServers_10_io_addressIn_ready),
    .io_addressIn_valid(casServers_10_io_addressIn_valid),
    .io_addressIn_bits(casServers_10_io_addressIn_bits),
    .io_addressOut_ready(casServers_10_io_addressOut_ready),
    .io_addressOut_valid(casServers_10_io_addressOut_valid),
    .io_addressOut_bits(casServers_10_io_addressOut_bits)
  );
  contAddrServer casServers_11 ( // @[contNetwork.scala 17:53]
    .clock(casServers_11_clock),
    .reset(casServers_11_reset),
    .io_addressIn_ready(casServers_11_io_addressIn_ready),
    .io_addressIn_valid(casServers_11_io_addressIn_valid),
    .io_addressIn_bits(casServers_11_io_addressIn_bits),
    .io_addressOut_ready(casServers_11_io_addressOut_ready),
    .io_addressOut_valid(casServers_11_io_addressOut_valid),
    .io_addressOut_bits(casServers_11_io_addressOut_bits)
  );
  contAddrServer casServers_12 ( // @[contNetwork.scala 17:53]
    .clock(casServers_12_clock),
    .reset(casServers_12_reset),
    .io_addressIn_ready(casServers_12_io_addressIn_ready),
    .io_addressIn_valid(casServers_12_io_addressIn_valid),
    .io_addressIn_bits(casServers_12_io_addressIn_bits),
    .io_addressOut_ready(casServers_12_io_addressOut_ready),
    .io_addressOut_valid(casServers_12_io_addressOut_valid),
    .io_addressOut_bits(casServers_12_io_addressOut_bits)
  );
  contAddrServer casServers_13 ( // @[contNetwork.scala 17:53]
    .clock(casServers_13_clock),
    .reset(casServers_13_reset),
    .io_addressIn_ready(casServers_13_io_addressIn_ready),
    .io_addressIn_valid(casServers_13_io_addressIn_valid),
    .io_addressIn_bits(casServers_13_io_addressIn_bits),
    .io_addressOut_ready(casServers_13_io_addressOut_ready),
    .io_addressOut_valid(casServers_13_io_addressOut_valid),
    .io_addressOut_bits(casServers_13_io_addressOut_bits)
  );
  contAddrServer casServers_14 ( // @[contNetwork.scala 17:53]
    .clock(casServers_14_clock),
    .reset(casServers_14_reset),
    .io_addressIn_ready(casServers_14_io_addressIn_ready),
    .io_addressIn_valid(casServers_14_io_addressIn_valid),
    .io_addressIn_bits(casServers_14_io_addressIn_bits),
    .io_addressOut_ready(casServers_14_io_addressOut_ready),
    .io_addressOut_valid(casServers_14_io_addressOut_valid),
    .io_addressOut_bits(casServers_14_io_addressOut_bits)
  );
  contAddrServer casServers_15 ( // @[contNetwork.scala 17:53]
    .clock(casServers_15_clock),
    .reset(casServers_15_reset),
    .io_addressIn_ready(casServers_15_io_addressIn_ready),
    .io_addressIn_valid(casServers_15_io_addressIn_valid),
    .io_addressIn_bits(casServers_15_io_addressIn_bits),
    .io_addressOut_ready(casServers_15_io_addressOut_ready),
    .io_addressOut_valid(casServers_15_io_addressOut_valid),
    .io_addressOut_bits(casServers_15_io_addressOut_bits)
  );
  contAddrServer casServers_16 ( // @[contNetwork.scala 17:53]
    .clock(casServers_16_clock),
    .reset(casServers_16_reset),
    .io_addressIn_ready(casServers_16_io_addressIn_ready),
    .io_addressIn_valid(casServers_16_io_addressIn_valid),
    .io_addressIn_bits(casServers_16_io_addressIn_bits),
    .io_addressOut_ready(casServers_16_io_addressOut_ready),
    .io_addressOut_valid(casServers_16_io_addressOut_valid),
    .io_addressOut_bits(casServers_16_io_addressOut_bits)
  );
  contAddrServer casServers_17 ( // @[contNetwork.scala 17:53]
    .clock(casServers_17_clock),
    .reset(casServers_17_reset),
    .io_addressIn_ready(casServers_17_io_addressIn_ready),
    .io_addressIn_valid(casServers_17_io_addressIn_valid),
    .io_addressIn_bits(casServers_17_io_addressIn_bits),
    .io_addressOut_ready(casServers_17_io_addressOut_ready),
    .io_addressOut_valid(casServers_17_io_addressOut_valid),
    .io_addressOut_bits(casServers_17_io_addressOut_bits)
  );
  contAddrServer casServers_18 ( // @[contNetwork.scala 17:53]
    .clock(casServers_18_clock),
    .reset(casServers_18_reset),
    .io_addressIn_ready(casServers_18_io_addressIn_ready),
    .io_addressIn_valid(casServers_18_io_addressIn_valid),
    .io_addressIn_bits(casServers_18_io_addressIn_bits),
    .io_addressOut_ready(casServers_18_io_addressOut_ready),
    .io_addressOut_valid(casServers_18_io_addressOut_valid),
    .io_addressOut_bits(casServers_18_io_addressOut_bits)
  );
  contAddrServer casServers_19 ( // @[contNetwork.scala 17:53]
    .clock(casServers_19_clock),
    .reset(casServers_19_reset),
    .io_addressIn_ready(casServers_19_io_addressIn_ready),
    .io_addressIn_valid(casServers_19_io_addressIn_valid),
    .io_addressIn_bits(casServers_19_io_addressIn_bits),
    .io_addressOut_ready(casServers_19_io_addressOut_ready),
    .io_addressOut_valid(casServers_19_io_addressOut_valid),
    .io_addressOut_bits(casServers_19_io_addressOut_bits)
  );
  contAddrServer casServers_20 ( // @[contNetwork.scala 17:53]
    .clock(casServers_20_clock),
    .reset(casServers_20_reset),
    .io_addressIn_ready(casServers_20_io_addressIn_ready),
    .io_addressIn_valid(casServers_20_io_addressIn_valid),
    .io_addressIn_bits(casServers_20_io_addressIn_bits),
    .io_addressOut_ready(casServers_20_io_addressOut_ready),
    .io_addressOut_valid(casServers_20_io_addressOut_valid),
    .io_addressOut_bits(casServers_20_io_addressOut_bits)
  );
  contAddrServer casServers_21 ( // @[contNetwork.scala 17:53]
    .clock(casServers_21_clock),
    .reset(casServers_21_reset),
    .io_addressIn_ready(casServers_21_io_addressIn_ready),
    .io_addressIn_valid(casServers_21_io_addressIn_valid),
    .io_addressIn_bits(casServers_21_io_addressIn_bits),
    .io_addressOut_ready(casServers_21_io_addressOut_ready),
    .io_addressOut_valid(casServers_21_io_addressOut_valid),
    .io_addressOut_bits(casServers_21_io_addressOut_bits)
  );
  contAddrServer casServers_22 ( // @[contNetwork.scala 17:53]
    .clock(casServers_22_clock),
    .reset(casServers_22_reset),
    .io_addressIn_ready(casServers_22_io_addressIn_ready),
    .io_addressIn_valid(casServers_22_io_addressIn_valid),
    .io_addressIn_bits(casServers_22_io_addressIn_bits),
    .io_addressOut_ready(casServers_22_io_addressOut_ready),
    .io_addressOut_valid(casServers_22_io_addressOut_valid),
    .io_addressOut_bits(casServers_22_io_addressOut_bits)
  );
  contAddrServer casServers_23 ( // @[contNetwork.scala 17:53]
    .clock(casServers_23_clock),
    .reset(casServers_23_reset),
    .io_addressIn_ready(casServers_23_io_addressIn_ready),
    .io_addressIn_valid(casServers_23_io_addressIn_valid),
    .io_addressIn_bits(casServers_23_io_addressIn_bits),
    .io_addressOut_ready(casServers_23_io_addressOut_ready),
    .io_addressOut_valid(casServers_23_io_addressOut_valid),
    .io_addressOut_bits(casServers_23_io_addressOut_bits)
  );
  contAddrServer casServers_24 ( // @[contNetwork.scala 17:53]
    .clock(casServers_24_clock),
    .reset(casServers_24_reset),
    .io_addressIn_ready(casServers_24_io_addressIn_ready),
    .io_addressIn_valid(casServers_24_io_addressIn_valid),
    .io_addressIn_bits(casServers_24_io_addressIn_bits),
    .io_addressOut_ready(casServers_24_io_addressOut_ready),
    .io_addressOut_valid(casServers_24_io_addressOut_valid),
    .io_addressOut_bits(casServers_24_io_addressOut_bits)
  );
  contAddrServer casServers_25 ( // @[contNetwork.scala 17:53]
    .clock(casServers_25_clock),
    .reset(casServers_25_reset),
    .io_addressIn_ready(casServers_25_io_addressIn_ready),
    .io_addressIn_valid(casServers_25_io_addressIn_valid),
    .io_addressIn_bits(casServers_25_io_addressIn_bits),
    .io_addressOut_ready(casServers_25_io_addressOut_ready),
    .io_addressOut_valid(casServers_25_io_addressOut_valid),
    .io_addressOut_bits(casServers_25_io_addressOut_bits)
  );
  contAddrServer casServers_26 ( // @[contNetwork.scala 17:53]
    .clock(casServers_26_clock),
    .reset(casServers_26_reset),
    .io_addressIn_ready(casServers_26_io_addressIn_ready),
    .io_addressIn_valid(casServers_26_io_addressIn_valid),
    .io_addressIn_bits(casServers_26_io_addressIn_bits),
    .io_addressOut_ready(casServers_26_io_addressOut_ready),
    .io_addressOut_valid(casServers_26_io_addressOut_valid),
    .io_addressOut_bits(casServers_26_io_addressOut_bits)
  );
  contAddrServer casServers_27 ( // @[contNetwork.scala 17:53]
    .clock(casServers_27_clock),
    .reset(casServers_27_reset),
    .io_addressIn_ready(casServers_27_io_addressIn_ready),
    .io_addressIn_valid(casServers_27_io_addressIn_valid),
    .io_addressIn_bits(casServers_27_io_addressIn_bits),
    .io_addressOut_ready(casServers_27_io_addressOut_ready),
    .io_addressOut_valid(casServers_27_io_addressOut_valid),
    .io_addressOut_bits(casServers_27_io_addressOut_bits)
  );
  contAddrServer casServers_28 ( // @[contNetwork.scala 17:53]
    .clock(casServers_28_clock),
    .reset(casServers_28_reset),
    .io_addressIn_ready(casServers_28_io_addressIn_ready),
    .io_addressIn_valid(casServers_28_io_addressIn_valid),
    .io_addressIn_bits(casServers_28_io_addressIn_bits),
    .io_addressOut_ready(casServers_28_io_addressOut_ready),
    .io_addressOut_valid(casServers_28_io_addressOut_valid),
    .io_addressOut_bits(casServers_28_io_addressOut_bits)
  );
  contAddrServer casServers_29 ( // @[contNetwork.scala 17:53]
    .clock(casServers_29_clock),
    .reset(casServers_29_reset),
    .io_addressIn_ready(casServers_29_io_addressIn_ready),
    .io_addressIn_valid(casServers_29_io_addressIn_valid),
    .io_addressIn_bits(casServers_29_io_addressIn_bits),
    .io_addressOut_ready(casServers_29_io_addressOut_ready),
    .io_addressOut_valid(casServers_29_io_addressOut_valid),
    .io_addressOut_bits(casServers_29_io_addressOut_bits)
  );
  contAddrServer casServers_30 ( // @[contNetwork.scala 17:53]
    .clock(casServers_30_clock),
    .reset(casServers_30_reset),
    .io_addressIn_ready(casServers_30_io_addressIn_ready),
    .io_addressIn_valid(casServers_30_io_addressIn_valid),
    .io_addressIn_bits(casServers_30_io_addressIn_bits),
    .io_addressOut_ready(casServers_30_io_addressOut_ready),
    .io_addressOut_valid(casServers_30_io_addressOut_valid),
    .io_addressOut_bits(casServers_30_io_addressOut_bits)
  );
  contAddrServer casServers_31 ( // @[contNetwork.scala 17:53]
    .clock(casServers_31_clock),
    .reset(casServers_31_reset),
    .io_addressIn_ready(casServers_31_io_addressIn_ready),
    .io_addressIn_valid(casServers_31_io_addressIn_valid),
    .io_addressIn_bits(casServers_31_io_addressIn_bits),
    .io_addressOut_ready(casServers_31_io_addressOut_ready),
    .io_addressOut_valid(casServers_31_io_addressOut_valid),
    .io_addressOut_bits(casServers_31_io_addressOut_bits)
  );
  contAddrServer casServers_32 ( // @[contNetwork.scala 17:53]
    .clock(casServers_32_clock),
    .reset(casServers_32_reset),
    .io_addressIn_ready(casServers_32_io_addressIn_ready),
    .io_addressIn_valid(casServers_32_io_addressIn_valid),
    .io_addressIn_bits(casServers_32_io_addressIn_bits),
    .io_addressOut_ready(casServers_32_io_addressOut_ready),
    .io_addressOut_valid(casServers_32_io_addressOut_valid),
    .io_addressOut_bits(casServers_32_io_addressOut_bits)
  );
  contAddrServer casServers_33 ( // @[contNetwork.scala 17:53]
    .clock(casServers_33_clock),
    .reset(casServers_33_reset),
    .io_addressIn_ready(casServers_33_io_addressIn_ready),
    .io_addressIn_valid(casServers_33_io_addressIn_valid),
    .io_addressIn_bits(casServers_33_io_addressIn_bits),
    .io_addressOut_ready(casServers_33_io_addressOut_ready),
    .io_addressOut_valid(casServers_33_io_addressOut_valid),
    .io_addressOut_bits(casServers_33_io_addressOut_bits)
  );
  contAddrServer casServers_34 ( // @[contNetwork.scala 17:53]
    .clock(casServers_34_clock),
    .reset(casServers_34_reset),
    .io_addressIn_ready(casServers_34_io_addressIn_ready),
    .io_addressIn_valid(casServers_34_io_addressIn_valid),
    .io_addressIn_bits(casServers_34_io_addressIn_bits),
    .io_addressOut_ready(casServers_34_io_addressOut_ready),
    .io_addressOut_valid(casServers_34_io_addressOut_valid),
    .io_addressOut_bits(casServers_34_io_addressOut_bits)
  );
  contAddrServer casServers_35 ( // @[contNetwork.scala 17:53]
    .clock(casServers_35_clock),
    .reset(casServers_35_reset),
    .io_addressIn_ready(casServers_35_io_addressIn_ready),
    .io_addressIn_valid(casServers_35_io_addressIn_valid),
    .io_addressIn_bits(casServers_35_io_addressIn_bits),
    .io_addressOut_ready(casServers_35_io_addressOut_ready),
    .io_addressOut_valid(casServers_35_io_addressOut_valid),
    .io_addressOut_bits(casServers_35_io_addressOut_bits)
  );
  contAddrServer casServers_36 ( // @[contNetwork.scala 17:53]
    .clock(casServers_36_clock),
    .reset(casServers_36_reset),
    .io_addressIn_ready(casServers_36_io_addressIn_ready),
    .io_addressIn_valid(casServers_36_io_addressIn_valid),
    .io_addressIn_bits(casServers_36_io_addressIn_bits),
    .io_addressOut_ready(casServers_36_io_addressOut_ready),
    .io_addressOut_valid(casServers_36_io_addressOut_valid),
    .io_addressOut_bits(casServers_36_io_addressOut_bits)
  );
  contAddrServer casServers_37 ( // @[contNetwork.scala 17:53]
    .clock(casServers_37_clock),
    .reset(casServers_37_reset),
    .io_addressIn_ready(casServers_37_io_addressIn_ready),
    .io_addressIn_valid(casServers_37_io_addressIn_valid),
    .io_addressIn_bits(casServers_37_io_addressIn_bits),
    .io_addressOut_ready(casServers_37_io_addressOut_ready),
    .io_addressOut_valid(casServers_37_io_addressOut_valid),
    .io_addressOut_bits(casServers_37_io_addressOut_bits)
  );
  contAddrServer casServers_38 ( // @[contNetwork.scala 17:53]
    .clock(casServers_38_clock),
    .reset(casServers_38_reset),
    .io_addressIn_ready(casServers_38_io_addressIn_ready),
    .io_addressIn_valid(casServers_38_io_addressIn_valid),
    .io_addressIn_bits(casServers_38_io_addressIn_bits),
    .io_addressOut_ready(casServers_38_io_addressOut_ready),
    .io_addressOut_valid(casServers_38_io_addressOut_valid),
    .io_addressOut_bits(casServers_38_io_addressOut_bits)
  );
  contAddrServer casServers_39 ( // @[contNetwork.scala 17:53]
    .clock(casServers_39_clock),
    .reset(casServers_39_reset),
    .io_addressIn_ready(casServers_39_io_addressIn_ready),
    .io_addressIn_valid(casServers_39_io_addressIn_valid),
    .io_addressIn_bits(casServers_39_io_addressIn_bits),
    .io_addressOut_ready(casServers_39_io_addressOut_ready),
    .io_addressOut_valid(casServers_39_io_addressOut_valid),
    .io_addressOut_bits(casServers_39_io_addressOut_bits)
  );
  contAddrServer casServers_40 ( // @[contNetwork.scala 17:53]
    .clock(casServers_40_clock),
    .reset(casServers_40_reset),
    .io_addressIn_ready(casServers_40_io_addressIn_ready),
    .io_addressIn_valid(casServers_40_io_addressIn_valid),
    .io_addressIn_bits(casServers_40_io_addressIn_bits),
    .io_addressOut_ready(casServers_40_io_addressOut_ready),
    .io_addressOut_valid(casServers_40_io_addressOut_valid),
    .io_addressOut_bits(casServers_40_io_addressOut_bits)
  );
  contAddrServer casServers_41 ( // @[contNetwork.scala 17:53]
    .clock(casServers_41_clock),
    .reset(casServers_41_reset),
    .io_addressIn_ready(casServers_41_io_addressIn_ready),
    .io_addressIn_valid(casServers_41_io_addressIn_valid),
    .io_addressIn_bits(casServers_41_io_addressIn_bits),
    .io_addressOut_ready(casServers_41_io_addressOut_ready),
    .io_addressOut_valid(casServers_41_io_addressOut_valid),
    .io_addressOut_bits(casServers_41_io_addressOut_bits)
  );
  contAddrServer casServers_42 ( // @[contNetwork.scala 17:53]
    .clock(casServers_42_clock),
    .reset(casServers_42_reset),
    .io_addressIn_ready(casServers_42_io_addressIn_ready),
    .io_addressIn_valid(casServers_42_io_addressIn_valid),
    .io_addressIn_bits(casServers_42_io_addressIn_bits),
    .io_addressOut_ready(casServers_42_io_addressOut_ready),
    .io_addressOut_valid(casServers_42_io_addressOut_valid),
    .io_addressOut_bits(casServers_42_io_addressOut_bits)
  );
  contAddrServer casServers_43 ( // @[contNetwork.scala 17:53]
    .clock(casServers_43_clock),
    .reset(casServers_43_reset),
    .io_addressIn_ready(casServers_43_io_addressIn_ready),
    .io_addressIn_valid(casServers_43_io_addressIn_valid),
    .io_addressIn_bits(casServers_43_io_addressIn_bits),
    .io_addressOut_ready(casServers_43_io_addressOut_ready),
    .io_addressOut_valid(casServers_43_io_addressOut_valid),
    .io_addressOut_bits(casServers_43_io_addressOut_bits)
  );
  contAddrServer casServers_44 ( // @[contNetwork.scala 17:53]
    .clock(casServers_44_clock),
    .reset(casServers_44_reset),
    .io_addressIn_ready(casServers_44_io_addressIn_ready),
    .io_addressIn_valid(casServers_44_io_addressIn_valid),
    .io_addressIn_bits(casServers_44_io_addressIn_bits),
    .io_addressOut_ready(casServers_44_io_addressOut_ready),
    .io_addressOut_valid(casServers_44_io_addressOut_valid),
    .io_addressOut_bits(casServers_44_io_addressOut_bits)
  );
  contAddrServer casServers_45 ( // @[contNetwork.scala 17:53]
    .clock(casServers_45_clock),
    .reset(casServers_45_reset),
    .io_addressIn_ready(casServers_45_io_addressIn_ready),
    .io_addressIn_valid(casServers_45_io_addressIn_valid),
    .io_addressIn_bits(casServers_45_io_addressIn_bits),
    .io_addressOut_ready(casServers_45_io_addressOut_ready),
    .io_addressOut_valid(casServers_45_io_addressOut_valid),
    .io_addressOut_bits(casServers_45_io_addressOut_bits)
  );
  contAddrServer casServers_46 ( // @[contNetwork.scala 17:53]
    .clock(casServers_46_clock),
    .reset(casServers_46_reset),
    .io_addressIn_ready(casServers_46_io_addressIn_ready),
    .io_addressIn_valid(casServers_46_io_addressIn_valid),
    .io_addressIn_bits(casServers_46_io_addressIn_bits),
    .io_addressOut_ready(casServers_46_io_addressOut_ready),
    .io_addressOut_valid(casServers_46_io_addressOut_valid),
    .io_addressOut_bits(casServers_46_io_addressOut_bits)
  );
  contAddrServer casServers_47 ( // @[contNetwork.scala 17:53]
    .clock(casServers_47_clock),
    .reset(casServers_47_reset),
    .io_addressIn_ready(casServers_47_io_addressIn_ready),
    .io_addressIn_valid(casServers_47_io_addressIn_valid),
    .io_addressIn_bits(casServers_47_io_addressIn_bits),
    .io_addressOut_ready(casServers_47_io_addressOut_ready),
    .io_addressOut_valid(casServers_47_io_addressOut_valid),
    .io_addressOut_bits(casServers_47_io_addressOut_bits)
  );
  contAddrServer casServers_48 ( // @[contNetwork.scala 17:53]
    .clock(casServers_48_clock),
    .reset(casServers_48_reset),
    .io_addressIn_ready(casServers_48_io_addressIn_ready),
    .io_addressIn_valid(casServers_48_io_addressIn_valid),
    .io_addressIn_bits(casServers_48_io_addressIn_bits),
    .io_addressOut_ready(casServers_48_io_addressOut_ready),
    .io_addressOut_valid(casServers_48_io_addressOut_valid),
    .io_addressOut_bits(casServers_48_io_addressOut_bits)
  );
  contAddrServer casServers_49 ( // @[contNetwork.scala 17:53]
    .clock(casServers_49_clock),
    .reset(casServers_49_reset),
    .io_addressIn_ready(casServers_49_io_addressIn_ready),
    .io_addressIn_valid(casServers_49_io_addressIn_valid),
    .io_addressIn_bits(casServers_49_io_addressIn_bits),
    .io_addressOut_ready(casServers_49_io_addressOut_ready),
    .io_addressOut_valid(casServers_49_io_addressOut_valid),
    .io_addressOut_bits(casServers_49_io_addressOut_bits)
  );
  contAddrServer casServers_50 ( // @[contNetwork.scala 17:53]
    .clock(casServers_50_clock),
    .reset(casServers_50_reset),
    .io_addressIn_ready(casServers_50_io_addressIn_ready),
    .io_addressIn_valid(casServers_50_io_addressIn_valid),
    .io_addressIn_bits(casServers_50_io_addressIn_bits),
    .io_addressOut_ready(casServers_50_io_addressOut_ready),
    .io_addressOut_valid(casServers_50_io_addressOut_valid),
    .io_addressOut_bits(casServers_50_io_addressOut_bits)
  );
  contAddrServer casServers_51 ( // @[contNetwork.scala 17:53]
    .clock(casServers_51_clock),
    .reset(casServers_51_reset),
    .io_addressIn_ready(casServers_51_io_addressIn_ready),
    .io_addressIn_valid(casServers_51_io_addressIn_valid),
    .io_addressIn_bits(casServers_51_io_addressIn_bits),
    .io_addressOut_ready(casServers_51_io_addressOut_ready),
    .io_addressOut_valid(casServers_51_io_addressOut_valid),
    .io_addressOut_bits(casServers_51_io_addressOut_bits)
  );
  contAddrServer casServers_52 ( // @[contNetwork.scala 17:53]
    .clock(casServers_52_clock),
    .reset(casServers_52_reset),
    .io_addressIn_ready(casServers_52_io_addressIn_ready),
    .io_addressIn_valid(casServers_52_io_addressIn_valid),
    .io_addressIn_bits(casServers_52_io_addressIn_bits),
    .io_addressOut_ready(casServers_52_io_addressOut_ready),
    .io_addressOut_valid(casServers_52_io_addressOut_valid),
    .io_addressOut_bits(casServers_52_io_addressOut_bits)
  );
  contAddrServer casServers_53 ( // @[contNetwork.scala 17:53]
    .clock(casServers_53_clock),
    .reset(casServers_53_reset),
    .io_addressIn_ready(casServers_53_io_addressIn_ready),
    .io_addressIn_valid(casServers_53_io_addressIn_valid),
    .io_addressIn_bits(casServers_53_io_addressIn_bits),
    .io_addressOut_ready(casServers_53_io_addressOut_ready),
    .io_addressOut_valid(casServers_53_io_addressOut_valid),
    .io_addressOut_bits(casServers_53_io_addressOut_bits)
  );
  contAddrServer casServers_54 ( // @[contNetwork.scala 17:53]
    .clock(casServers_54_clock),
    .reset(casServers_54_reset),
    .io_addressIn_ready(casServers_54_io_addressIn_ready),
    .io_addressIn_valid(casServers_54_io_addressIn_valid),
    .io_addressIn_bits(casServers_54_io_addressIn_bits),
    .io_addressOut_ready(casServers_54_io_addressOut_ready),
    .io_addressOut_valid(casServers_54_io_addressOut_valid),
    .io_addressOut_bits(casServers_54_io_addressOut_bits)
  );
  contAddrServer casServers_55 ( // @[contNetwork.scala 17:53]
    .clock(casServers_55_clock),
    .reset(casServers_55_reset),
    .io_addressIn_ready(casServers_55_io_addressIn_ready),
    .io_addressIn_valid(casServers_55_io_addressIn_valid),
    .io_addressIn_bits(casServers_55_io_addressIn_bits),
    .io_addressOut_ready(casServers_55_io_addressOut_ready),
    .io_addressOut_valid(casServers_55_io_addressOut_valid),
    .io_addressOut_bits(casServers_55_io_addressOut_bits)
  );
  contAddrServer casServers_56 ( // @[contNetwork.scala 17:53]
    .clock(casServers_56_clock),
    .reset(casServers_56_reset),
    .io_addressIn_ready(casServers_56_io_addressIn_ready),
    .io_addressIn_valid(casServers_56_io_addressIn_valid),
    .io_addressIn_bits(casServers_56_io_addressIn_bits),
    .io_addressOut_ready(casServers_56_io_addressOut_ready),
    .io_addressOut_valid(casServers_56_io_addressOut_valid),
    .io_addressOut_bits(casServers_56_io_addressOut_bits)
  );
  contAddrServer casServers_57 ( // @[contNetwork.scala 17:53]
    .clock(casServers_57_clock),
    .reset(casServers_57_reset),
    .io_addressIn_ready(casServers_57_io_addressIn_ready),
    .io_addressIn_valid(casServers_57_io_addressIn_valid),
    .io_addressIn_bits(casServers_57_io_addressIn_bits),
    .io_addressOut_ready(casServers_57_io_addressOut_ready),
    .io_addressOut_valid(casServers_57_io_addressOut_valid),
    .io_addressOut_bits(casServers_57_io_addressOut_bits)
  );
  contAddrServer casServers_58 ( // @[contNetwork.scala 17:53]
    .clock(casServers_58_clock),
    .reset(casServers_58_reset),
    .io_addressIn_ready(casServers_58_io_addressIn_ready),
    .io_addressIn_valid(casServers_58_io_addressIn_valid),
    .io_addressIn_bits(casServers_58_io_addressIn_bits),
    .io_addressOut_ready(casServers_58_io_addressOut_ready),
    .io_addressOut_valid(casServers_58_io_addressOut_valid),
    .io_addressOut_bits(casServers_58_io_addressOut_bits)
  );
  contAddrServer casServers_59 ( // @[contNetwork.scala 17:53]
    .clock(casServers_59_clock),
    .reset(casServers_59_reset),
    .io_addressIn_ready(casServers_59_io_addressIn_ready),
    .io_addressIn_valid(casServers_59_io_addressIn_valid),
    .io_addressIn_bits(casServers_59_io_addressIn_bits),
    .io_addressOut_ready(casServers_59_io_addressOut_ready),
    .io_addressOut_valid(casServers_59_io_addressOut_valid),
    .io_addressOut_bits(casServers_59_io_addressOut_bits)
  );
  contAddrServer casServers_60 ( // @[contNetwork.scala 17:53]
    .clock(casServers_60_clock),
    .reset(casServers_60_reset),
    .io_addressIn_ready(casServers_60_io_addressIn_ready),
    .io_addressIn_valid(casServers_60_io_addressIn_valid),
    .io_addressIn_bits(casServers_60_io_addressIn_bits),
    .io_addressOut_ready(casServers_60_io_addressOut_ready),
    .io_addressOut_valid(casServers_60_io_addressOut_valid),
    .io_addressOut_bits(casServers_60_io_addressOut_bits)
  );
  contAddrServer casServers_61 ( // @[contNetwork.scala 17:53]
    .clock(casServers_61_clock),
    .reset(casServers_61_reset),
    .io_addressIn_ready(casServers_61_io_addressIn_ready),
    .io_addressIn_valid(casServers_61_io_addressIn_valid),
    .io_addressIn_bits(casServers_61_io_addressIn_bits),
    .io_addressOut_ready(casServers_61_io_addressOut_ready),
    .io_addressOut_valid(casServers_61_io_addressOut_valid),
    .io_addressOut_bits(casServers_61_io_addressOut_bits)
  );
  contAddrServer casServers_62 ( // @[contNetwork.scala 17:53]
    .clock(casServers_62_clock),
    .reset(casServers_62_reset),
    .io_addressIn_ready(casServers_62_io_addressIn_ready),
    .io_addressIn_valid(casServers_62_io_addressIn_valid),
    .io_addressIn_bits(casServers_62_io_addressIn_bits),
    .io_addressOut_ready(casServers_62_io_addressOut_ready),
    .io_addressOut_valid(casServers_62_io_addressOut_valid),
    .io_addressOut_bits(casServers_62_io_addressOut_bits)
  );
  contAddrServer casServers_63 ( // @[contNetwork.scala 17:53]
    .clock(casServers_63_clock),
    .reset(casServers_63_reset),
    .io_addressIn_ready(casServers_63_io_addressIn_ready),
    .io_addressIn_valid(casServers_63_io_addressIn_valid),
    .io_addressIn_bits(casServers_63_io_addressIn_bits),
    .io_addressOut_ready(casServers_63_io_addressOut_ready),
    .io_addressOut_valid(casServers_63_io_addressOut_valid),
    .io_addressOut_bits(casServers_63_io_addressOut_bits)
  );
  contQueue queues_0 ( // @[contNetwork.scala 18:53]
    .clock(queues_0_clock),
    .reset(queues_0_reset),
    .io_addressIn_ready(queues_0_io_addressIn_ready),
    .io_addressIn_valid(queues_0_io_addressIn_valid),
    .io_addressIn_bits(queues_0_io_addressIn_bits),
    .io_addressOut_ready(queues_0_io_addressOut_ready),
    .io_addressOut_valid(queues_0_io_addressOut_valid),
    .io_addressOut_bits(queues_0_io_addressOut_bits)
  );
  contQueue queues_1 ( // @[contNetwork.scala 18:53]
    .clock(queues_1_clock),
    .reset(queues_1_reset),
    .io_addressIn_ready(queues_1_io_addressIn_ready),
    .io_addressIn_valid(queues_1_io_addressIn_valid),
    .io_addressIn_bits(queues_1_io_addressIn_bits),
    .io_addressOut_ready(queues_1_io_addressOut_ready),
    .io_addressOut_valid(queues_1_io_addressOut_valid),
    .io_addressOut_bits(queues_1_io_addressOut_bits)
  );
  contQueue queues_2 ( // @[contNetwork.scala 18:53]
    .clock(queues_2_clock),
    .reset(queues_2_reset),
    .io_addressIn_ready(queues_2_io_addressIn_ready),
    .io_addressIn_valid(queues_2_io_addressIn_valid),
    .io_addressIn_bits(queues_2_io_addressIn_bits),
    .io_addressOut_ready(queues_2_io_addressOut_ready),
    .io_addressOut_valid(queues_2_io_addressOut_valid),
    .io_addressOut_bits(queues_2_io_addressOut_bits)
  );
  contQueue queues_3 ( // @[contNetwork.scala 18:53]
    .clock(queues_3_clock),
    .reset(queues_3_reset),
    .io_addressIn_ready(queues_3_io_addressIn_ready),
    .io_addressIn_valid(queues_3_io_addressIn_valid),
    .io_addressIn_bits(queues_3_io_addressIn_bits),
    .io_addressOut_ready(queues_3_io_addressOut_ready),
    .io_addressOut_valid(queues_3_io_addressOut_valid),
    .io_addressOut_bits(queues_3_io_addressOut_bits)
  );
  contQueue queues_4 ( // @[contNetwork.scala 18:53]
    .clock(queues_4_clock),
    .reset(queues_4_reset),
    .io_addressIn_ready(queues_4_io_addressIn_ready),
    .io_addressIn_valid(queues_4_io_addressIn_valid),
    .io_addressIn_bits(queues_4_io_addressIn_bits),
    .io_addressOut_ready(queues_4_io_addressOut_ready),
    .io_addressOut_valid(queues_4_io_addressOut_valid),
    .io_addressOut_bits(queues_4_io_addressOut_bits)
  );
  contQueue queues_5 ( // @[contNetwork.scala 18:53]
    .clock(queues_5_clock),
    .reset(queues_5_reset),
    .io_addressIn_ready(queues_5_io_addressIn_ready),
    .io_addressIn_valid(queues_5_io_addressIn_valid),
    .io_addressIn_bits(queues_5_io_addressIn_bits),
    .io_addressOut_ready(queues_5_io_addressOut_ready),
    .io_addressOut_valid(queues_5_io_addressOut_valid),
    .io_addressOut_bits(queues_5_io_addressOut_bits)
  );
  contQueue queues_6 ( // @[contNetwork.scala 18:53]
    .clock(queues_6_clock),
    .reset(queues_6_reset),
    .io_addressIn_ready(queues_6_io_addressIn_ready),
    .io_addressIn_valid(queues_6_io_addressIn_valid),
    .io_addressIn_bits(queues_6_io_addressIn_bits),
    .io_addressOut_ready(queues_6_io_addressOut_ready),
    .io_addressOut_valid(queues_6_io_addressOut_valid),
    .io_addressOut_bits(queues_6_io_addressOut_bits)
  );
  contQueue queues_7 ( // @[contNetwork.scala 18:53]
    .clock(queues_7_clock),
    .reset(queues_7_reset),
    .io_addressIn_ready(queues_7_io_addressIn_ready),
    .io_addressIn_valid(queues_7_io_addressIn_valid),
    .io_addressIn_bits(queues_7_io_addressIn_bits),
    .io_addressOut_ready(queues_7_io_addressOut_ready),
    .io_addressOut_valid(queues_7_io_addressOut_valid),
    .io_addressOut_bits(queues_7_io_addressOut_bits)
  );
  contQueue queues_8 ( // @[contNetwork.scala 18:53]
    .clock(queues_8_clock),
    .reset(queues_8_reset),
    .io_addressIn_ready(queues_8_io_addressIn_ready),
    .io_addressIn_valid(queues_8_io_addressIn_valid),
    .io_addressIn_bits(queues_8_io_addressIn_bits),
    .io_addressOut_ready(queues_8_io_addressOut_ready),
    .io_addressOut_valid(queues_8_io_addressOut_valid),
    .io_addressOut_bits(queues_8_io_addressOut_bits)
  );
  contQueue queues_9 ( // @[contNetwork.scala 18:53]
    .clock(queues_9_clock),
    .reset(queues_9_reset),
    .io_addressIn_ready(queues_9_io_addressIn_ready),
    .io_addressIn_valid(queues_9_io_addressIn_valid),
    .io_addressIn_bits(queues_9_io_addressIn_bits),
    .io_addressOut_ready(queues_9_io_addressOut_ready),
    .io_addressOut_valid(queues_9_io_addressOut_valid),
    .io_addressOut_bits(queues_9_io_addressOut_bits)
  );
  contQueue queues_10 ( // @[contNetwork.scala 18:53]
    .clock(queues_10_clock),
    .reset(queues_10_reset),
    .io_addressIn_ready(queues_10_io_addressIn_ready),
    .io_addressIn_valid(queues_10_io_addressIn_valid),
    .io_addressIn_bits(queues_10_io_addressIn_bits),
    .io_addressOut_ready(queues_10_io_addressOut_ready),
    .io_addressOut_valid(queues_10_io_addressOut_valid),
    .io_addressOut_bits(queues_10_io_addressOut_bits)
  );
  contQueue queues_11 ( // @[contNetwork.scala 18:53]
    .clock(queues_11_clock),
    .reset(queues_11_reset),
    .io_addressIn_ready(queues_11_io_addressIn_ready),
    .io_addressIn_valid(queues_11_io_addressIn_valid),
    .io_addressIn_bits(queues_11_io_addressIn_bits),
    .io_addressOut_ready(queues_11_io_addressOut_ready),
    .io_addressOut_valid(queues_11_io_addressOut_valid),
    .io_addressOut_bits(queues_11_io_addressOut_bits)
  );
  contQueue queues_12 ( // @[contNetwork.scala 18:53]
    .clock(queues_12_clock),
    .reset(queues_12_reset),
    .io_addressIn_ready(queues_12_io_addressIn_ready),
    .io_addressIn_valid(queues_12_io_addressIn_valid),
    .io_addressIn_bits(queues_12_io_addressIn_bits),
    .io_addressOut_ready(queues_12_io_addressOut_ready),
    .io_addressOut_valid(queues_12_io_addressOut_valid),
    .io_addressOut_bits(queues_12_io_addressOut_bits)
  );
  contQueue queues_13 ( // @[contNetwork.scala 18:53]
    .clock(queues_13_clock),
    .reset(queues_13_reset),
    .io_addressIn_ready(queues_13_io_addressIn_ready),
    .io_addressIn_valid(queues_13_io_addressIn_valid),
    .io_addressIn_bits(queues_13_io_addressIn_bits),
    .io_addressOut_ready(queues_13_io_addressOut_ready),
    .io_addressOut_valid(queues_13_io_addressOut_valid),
    .io_addressOut_bits(queues_13_io_addressOut_bits)
  );
  contQueue queues_14 ( // @[contNetwork.scala 18:53]
    .clock(queues_14_clock),
    .reset(queues_14_reset),
    .io_addressIn_ready(queues_14_io_addressIn_ready),
    .io_addressIn_valid(queues_14_io_addressIn_valid),
    .io_addressIn_bits(queues_14_io_addressIn_bits),
    .io_addressOut_ready(queues_14_io_addressOut_ready),
    .io_addressOut_valid(queues_14_io_addressOut_valid),
    .io_addressOut_bits(queues_14_io_addressOut_bits)
  );
  contQueue queues_15 ( // @[contNetwork.scala 18:53]
    .clock(queues_15_clock),
    .reset(queues_15_reset),
    .io_addressIn_ready(queues_15_io_addressIn_ready),
    .io_addressIn_valid(queues_15_io_addressIn_valid),
    .io_addressIn_bits(queues_15_io_addressIn_bits),
    .io_addressOut_ready(queues_15_io_addressOut_ready),
    .io_addressOut_valid(queues_15_io_addressOut_valid),
    .io_addressOut_bits(queues_15_io_addressOut_bits)
  );
  contQueue queues_16 ( // @[contNetwork.scala 18:53]
    .clock(queues_16_clock),
    .reset(queues_16_reset),
    .io_addressIn_ready(queues_16_io_addressIn_ready),
    .io_addressIn_valid(queues_16_io_addressIn_valid),
    .io_addressIn_bits(queues_16_io_addressIn_bits),
    .io_addressOut_ready(queues_16_io_addressOut_ready),
    .io_addressOut_valid(queues_16_io_addressOut_valid),
    .io_addressOut_bits(queues_16_io_addressOut_bits)
  );
  contQueue queues_17 ( // @[contNetwork.scala 18:53]
    .clock(queues_17_clock),
    .reset(queues_17_reset),
    .io_addressIn_ready(queues_17_io_addressIn_ready),
    .io_addressIn_valid(queues_17_io_addressIn_valid),
    .io_addressIn_bits(queues_17_io_addressIn_bits),
    .io_addressOut_ready(queues_17_io_addressOut_ready),
    .io_addressOut_valid(queues_17_io_addressOut_valid),
    .io_addressOut_bits(queues_17_io_addressOut_bits)
  );
  contQueue queues_18 ( // @[contNetwork.scala 18:53]
    .clock(queues_18_clock),
    .reset(queues_18_reset),
    .io_addressIn_ready(queues_18_io_addressIn_ready),
    .io_addressIn_valid(queues_18_io_addressIn_valid),
    .io_addressIn_bits(queues_18_io_addressIn_bits),
    .io_addressOut_ready(queues_18_io_addressOut_ready),
    .io_addressOut_valid(queues_18_io_addressOut_valid),
    .io_addressOut_bits(queues_18_io_addressOut_bits)
  );
  contQueue queues_19 ( // @[contNetwork.scala 18:53]
    .clock(queues_19_clock),
    .reset(queues_19_reset),
    .io_addressIn_ready(queues_19_io_addressIn_ready),
    .io_addressIn_valid(queues_19_io_addressIn_valid),
    .io_addressIn_bits(queues_19_io_addressIn_bits),
    .io_addressOut_ready(queues_19_io_addressOut_ready),
    .io_addressOut_valid(queues_19_io_addressOut_valid),
    .io_addressOut_bits(queues_19_io_addressOut_bits)
  );
  contQueue queues_20 ( // @[contNetwork.scala 18:53]
    .clock(queues_20_clock),
    .reset(queues_20_reset),
    .io_addressIn_ready(queues_20_io_addressIn_ready),
    .io_addressIn_valid(queues_20_io_addressIn_valid),
    .io_addressIn_bits(queues_20_io_addressIn_bits),
    .io_addressOut_ready(queues_20_io_addressOut_ready),
    .io_addressOut_valid(queues_20_io_addressOut_valid),
    .io_addressOut_bits(queues_20_io_addressOut_bits)
  );
  contQueue queues_21 ( // @[contNetwork.scala 18:53]
    .clock(queues_21_clock),
    .reset(queues_21_reset),
    .io_addressIn_ready(queues_21_io_addressIn_ready),
    .io_addressIn_valid(queues_21_io_addressIn_valid),
    .io_addressIn_bits(queues_21_io_addressIn_bits),
    .io_addressOut_ready(queues_21_io_addressOut_ready),
    .io_addressOut_valid(queues_21_io_addressOut_valid),
    .io_addressOut_bits(queues_21_io_addressOut_bits)
  );
  contQueue queues_22 ( // @[contNetwork.scala 18:53]
    .clock(queues_22_clock),
    .reset(queues_22_reset),
    .io_addressIn_ready(queues_22_io_addressIn_ready),
    .io_addressIn_valid(queues_22_io_addressIn_valid),
    .io_addressIn_bits(queues_22_io_addressIn_bits),
    .io_addressOut_ready(queues_22_io_addressOut_ready),
    .io_addressOut_valid(queues_22_io_addressOut_valid),
    .io_addressOut_bits(queues_22_io_addressOut_bits)
  );
  contQueue queues_23 ( // @[contNetwork.scala 18:53]
    .clock(queues_23_clock),
    .reset(queues_23_reset),
    .io_addressIn_ready(queues_23_io_addressIn_ready),
    .io_addressIn_valid(queues_23_io_addressIn_valid),
    .io_addressIn_bits(queues_23_io_addressIn_bits),
    .io_addressOut_ready(queues_23_io_addressOut_ready),
    .io_addressOut_valid(queues_23_io_addressOut_valid),
    .io_addressOut_bits(queues_23_io_addressOut_bits)
  );
  contQueue queues_24 ( // @[contNetwork.scala 18:53]
    .clock(queues_24_clock),
    .reset(queues_24_reset),
    .io_addressIn_ready(queues_24_io_addressIn_ready),
    .io_addressIn_valid(queues_24_io_addressIn_valid),
    .io_addressIn_bits(queues_24_io_addressIn_bits),
    .io_addressOut_ready(queues_24_io_addressOut_ready),
    .io_addressOut_valid(queues_24_io_addressOut_valid),
    .io_addressOut_bits(queues_24_io_addressOut_bits)
  );
  contQueue queues_25 ( // @[contNetwork.scala 18:53]
    .clock(queues_25_clock),
    .reset(queues_25_reset),
    .io_addressIn_ready(queues_25_io_addressIn_ready),
    .io_addressIn_valid(queues_25_io_addressIn_valid),
    .io_addressIn_bits(queues_25_io_addressIn_bits),
    .io_addressOut_ready(queues_25_io_addressOut_ready),
    .io_addressOut_valid(queues_25_io_addressOut_valid),
    .io_addressOut_bits(queues_25_io_addressOut_bits)
  );
  contQueue queues_26 ( // @[contNetwork.scala 18:53]
    .clock(queues_26_clock),
    .reset(queues_26_reset),
    .io_addressIn_ready(queues_26_io_addressIn_ready),
    .io_addressIn_valid(queues_26_io_addressIn_valid),
    .io_addressIn_bits(queues_26_io_addressIn_bits),
    .io_addressOut_ready(queues_26_io_addressOut_ready),
    .io_addressOut_valid(queues_26_io_addressOut_valid),
    .io_addressOut_bits(queues_26_io_addressOut_bits)
  );
  contQueue queues_27 ( // @[contNetwork.scala 18:53]
    .clock(queues_27_clock),
    .reset(queues_27_reset),
    .io_addressIn_ready(queues_27_io_addressIn_ready),
    .io_addressIn_valid(queues_27_io_addressIn_valid),
    .io_addressIn_bits(queues_27_io_addressIn_bits),
    .io_addressOut_ready(queues_27_io_addressOut_ready),
    .io_addressOut_valid(queues_27_io_addressOut_valid),
    .io_addressOut_bits(queues_27_io_addressOut_bits)
  );
  contQueue queues_28 ( // @[contNetwork.scala 18:53]
    .clock(queues_28_clock),
    .reset(queues_28_reset),
    .io_addressIn_ready(queues_28_io_addressIn_ready),
    .io_addressIn_valid(queues_28_io_addressIn_valid),
    .io_addressIn_bits(queues_28_io_addressIn_bits),
    .io_addressOut_ready(queues_28_io_addressOut_ready),
    .io_addressOut_valid(queues_28_io_addressOut_valid),
    .io_addressOut_bits(queues_28_io_addressOut_bits)
  );
  contQueue queues_29 ( // @[contNetwork.scala 18:53]
    .clock(queues_29_clock),
    .reset(queues_29_reset),
    .io_addressIn_ready(queues_29_io_addressIn_ready),
    .io_addressIn_valid(queues_29_io_addressIn_valid),
    .io_addressIn_bits(queues_29_io_addressIn_bits),
    .io_addressOut_ready(queues_29_io_addressOut_ready),
    .io_addressOut_valid(queues_29_io_addressOut_valid),
    .io_addressOut_bits(queues_29_io_addressOut_bits)
  );
  contQueue queues_30 ( // @[contNetwork.scala 18:53]
    .clock(queues_30_clock),
    .reset(queues_30_reset),
    .io_addressIn_ready(queues_30_io_addressIn_ready),
    .io_addressIn_valid(queues_30_io_addressIn_valid),
    .io_addressIn_bits(queues_30_io_addressIn_bits),
    .io_addressOut_ready(queues_30_io_addressOut_ready),
    .io_addressOut_valid(queues_30_io_addressOut_valid),
    .io_addressOut_bits(queues_30_io_addressOut_bits)
  );
  contQueue queues_31 ( // @[contNetwork.scala 18:53]
    .clock(queues_31_clock),
    .reset(queues_31_reset),
    .io_addressIn_ready(queues_31_io_addressIn_ready),
    .io_addressIn_valid(queues_31_io_addressIn_valid),
    .io_addressIn_bits(queues_31_io_addressIn_bits),
    .io_addressOut_ready(queues_31_io_addressOut_ready),
    .io_addressOut_valid(queues_31_io_addressOut_valid),
    .io_addressOut_bits(queues_31_io_addressOut_bits)
  );
  contQueue queues_32 ( // @[contNetwork.scala 18:53]
    .clock(queues_32_clock),
    .reset(queues_32_reset),
    .io_addressIn_ready(queues_32_io_addressIn_ready),
    .io_addressIn_valid(queues_32_io_addressIn_valid),
    .io_addressIn_bits(queues_32_io_addressIn_bits),
    .io_addressOut_ready(queues_32_io_addressOut_ready),
    .io_addressOut_valid(queues_32_io_addressOut_valid),
    .io_addressOut_bits(queues_32_io_addressOut_bits)
  );
  contQueue queues_33 ( // @[contNetwork.scala 18:53]
    .clock(queues_33_clock),
    .reset(queues_33_reset),
    .io_addressIn_ready(queues_33_io_addressIn_ready),
    .io_addressIn_valid(queues_33_io_addressIn_valid),
    .io_addressIn_bits(queues_33_io_addressIn_bits),
    .io_addressOut_ready(queues_33_io_addressOut_ready),
    .io_addressOut_valid(queues_33_io_addressOut_valid),
    .io_addressOut_bits(queues_33_io_addressOut_bits)
  );
  contQueue queues_34 ( // @[contNetwork.scala 18:53]
    .clock(queues_34_clock),
    .reset(queues_34_reset),
    .io_addressIn_ready(queues_34_io_addressIn_ready),
    .io_addressIn_valid(queues_34_io_addressIn_valid),
    .io_addressIn_bits(queues_34_io_addressIn_bits),
    .io_addressOut_ready(queues_34_io_addressOut_ready),
    .io_addressOut_valid(queues_34_io_addressOut_valid),
    .io_addressOut_bits(queues_34_io_addressOut_bits)
  );
  contQueue queues_35 ( // @[contNetwork.scala 18:53]
    .clock(queues_35_clock),
    .reset(queues_35_reset),
    .io_addressIn_ready(queues_35_io_addressIn_ready),
    .io_addressIn_valid(queues_35_io_addressIn_valid),
    .io_addressIn_bits(queues_35_io_addressIn_bits),
    .io_addressOut_ready(queues_35_io_addressOut_ready),
    .io_addressOut_valid(queues_35_io_addressOut_valid),
    .io_addressOut_bits(queues_35_io_addressOut_bits)
  );
  contQueue queues_36 ( // @[contNetwork.scala 18:53]
    .clock(queues_36_clock),
    .reset(queues_36_reset),
    .io_addressIn_ready(queues_36_io_addressIn_ready),
    .io_addressIn_valid(queues_36_io_addressIn_valid),
    .io_addressIn_bits(queues_36_io_addressIn_bits),
    .io_addressOut_ready(queues_36_io_addressOut_ready),
    .io_addressOut_valid(queues_36_io_addressOut_valid),
    .io_addressOut_bits(queues_36_io_addressOut_bits)
  );
  contQueue queues_37 ( // @[contNetwork.scala 18:53]
    .clock(queues_37_clock),
    .reset(queues_37_reset),
    .io_addressIn_ready(queues_37_io_addressIn_ready),
    .io_addressIn_valid(queues_37_io_addressIn_valid),
    .io_addressIn_bits(queues_37_io_addressIn_bits),
    .io_addressOut_ready(queues_37_io_addressOut_ready),
    .io_addressOut_valid(queues_37_io_addressOut_valid),
    .io_addressOut_bits(queues_37_io_addressOut_bits)
  );
  contQueue queues_38 ( // @[contNetwork.scala 18:53]
    .clock(queues_38_clock),
    .reset(queues_38_reset),
    .io_addressIn_ready(queues_38_io_addressIn_ready),
    .io_addressIn_valid(queues_38_io_addressIn_valid),
    .io_addressIn_bits(queues_38_io_addressIn_bits),
    .io_addressOut_ready(queues_38_io_addressOut_ready),
    .io_addressOut_valid(queues_38_io_addressOut_valid),
    .io_addressOut_bits(queues_38_io_addressOut_bits)
  );
  contQueue queues_39 ( // @[contNetwork.scala 18:53]
    .clock(queues_39_clock),
    .reset(queues_39_reset),
    .io_addressIn_ready(queues_39_io_addressIn_ready),
    .io_addressIn_valid(queues_39_io_addressIn_valid),
    .io_addressIn_bits(queues_39_io_addressIn_bits),
    .io_addressOut_ready(queues_39_io_addressOut_ready),
    .io_addressOut_valid(queues_39_io_addressOut_valid),
    .io_addressOut_bits(queues_39_io_addressOut_bits)
  );
  contQueue queues_40 ( // @[contNetwork.scala 18:53]
    .clock(queues_40_clock),
    .reset(queues_40_reset),
    .io_addressIn_ready(queues_40_io_addressIn_ready),
    .io_addressIn_valid(queues_40_io_addressIn_valid),
    .io_addressIn_bits(queues_40_io_addressIn_bits),
    .io_addressOut_ready(queues_40_io_addressOut_ready),
    .io_addressOut_valid(queues_40_io_addressOut_valid),
    .io_addressOut_bits(queues_40_io_addressOut_bits)
  );
  contQueue queues_41 ( // @[contNetwork.scala 18:53]
    .clock(queues_41_clock),
    .reset(queues_41_reset),
    .io_addressIn_ready(queues_41_io_addressIn_ready),
    .io_addressIn_valid(queues_41_io_addressIn_valid),
    .io_addressIn_bits(queues_41_io_addressIn_bits),
    .io_addressOut_ready(queues_41_io_addressOut_ready),
    .io_addressOut_valid(queues_41_io_addressOut_valid),
    .io_addressOut_bits(queues_41_io_addressOut_bits)
  );
  contQueue queues_42 ( // @[contNetwork.scala 18:53]
    .clock(queues_42_clock),
    .reset(queues_42_reset),
    .io_addressIn_ready(queues_42_io_addressIn_ready),
    .io_addressIn_valid(queues_42_io_addressIn_valid),
    .io_addressIn_bits(queues_42_io_addressIn_bits),
    .io_addressOut_ready(queues_42_io_addressOut_ready),
    .io_addressOut_valid(queues_42_io_addressOut_valid),
    .io_addressOut_bits(queues_42_io_addressOut_bits)
  );
  contQueue queues_43 ( // @[contNetwork.scala 18:53]
    .clock(queues_43_clock),
    .reset(queues_43_reset),
    .io_addressIn_ready(queues_43_io_addressIn_ready),
    .io_addressIn_valid(queues_43_io_addressIn_valid),
    .io_addressIn_bits(queues_43_io_addressIn_bits),
    .io_addressOut_ready(queues_43_io_addressOut_ready),
    .io_addressOut_valid(queues_43_io_addressOut_valid),
    .io_addressOut_bits(queues_43_io_addressOut_bits)
  );
  contQueue queues_44 ( // @[contNetwork.scala 18:53]
    .clock(queues_44_clock),
    .reset(queues_44_reset),
    .io_addressIn_ready(queues_44_io_addressIn_ready),
    .io_addressIn_valid(queues_44_io_addressIn_valid),
    .io_addressIn_bits(queues_44_io_addressIn_bits),
    .io_addressOut_ready(queues_44_io_addressOut_ready),
    .io_addressOut_valid(queues_44_io_addressOut_valid),
    .io_addressOut_bits(queues_44_io_addressOut_bits)
  );
  contQueue queues_45 ( // @[contNetwork.scala 18:53]
    .clock(queues_45_clock),
    .reset(queues_45_reset),
    .io_addressIn_ready(queues_45_io_addressIn_ready),
    .io_addressIn_valid(queues_45_io_addressIn_valid),
    .io_addressIn_bits(queues_45_io_addressIn_bits),
    .io_addressOut_ready(queues_45_io_addressOut_ready),
    .io_addressOut_valid(queues_45_io_addressOut_valid),
    .io_addressOut_bits(queues_45_io_addressOut_bits)
  );
  contQueue queues_46 ( // @[contNetwork.scala 18:53]
    .clock(queues_46_clock),
    .reset(queues_46_reset),
    .io_addressIn_ready(queues_46_io_addressIn_ready),
    .io_addressIn_valid(queues_46_io_addressIn_valid),
    .io_addressIn_bits(queues_46_io_addressIn_bits),
    .io_addressOut_ready(queues_46_io_addressOut_ready),
    .io_addressOut_valid(queues_46_io_addressOut_valid),
    .io_addressOut_bits(queues_46_io_addressOut_bits)
  );
  contQueue queues_47 ( // @[contNetwork.scala 18:53]
    .clock(queues_47_clock),
    .reset(queues_47_reset),
    .io_addressIn_ready(queues_47_io_addressIn_ready),
    .io_addressIn_valid(queues_47_io_addressIn_valid),
    .io_addressIn_bits(queues_47_io_addressIn_bits),
    .io_addressOut_ready(queues_47_io_addressOut_ready),
    .io_addressOut_valid(queues_47_io_addressOut_valid),
    .io_addressOut_bits(queues_47_io_addressOut_bits)
  );
  contQueue queues_48 ( // @[contNetwork.scala 18:53]
    .clock(queues_48_clock),
    .reset(queues_48_reset),
    .io_addressIn_ready(queues_48_io_addressIn_ready),
    .io_addressIn_valid(queues_48_io_addressIn_valid),
    .io_addressIn_bits(queues_48_io_addressIn_bits),
    .io_addressOut_ready(queues_48_io_addressOut_ready),
    .io_addressOut_valid(queues_48_io_addressOut_valid),
    .io_addressOut_bits(queues_48_io_addressOut_bits)
  );
  contQueue queues_49 ( // @[contNetwork.scala 18:53]
    .clock(queues_49_clock),
    .reset(queues_49_reset),
    .io_addressIn_ready(queues_49_io_addressIn_ready),
    .io_addressIn_valid(queues_49_io_addressIn_valid),
    .io_addressIn_bits(queues_49_io_addressIn_bits),
    .io_addressOut_ready(queues_49_io_addressOut_ready),
    .io_addressOut_valid(queues_49_io_addressOut_valid),
    .io_addressOut_bits(queues_49_io_addressOut_bits)
  );
  contQueue queues_50 ( // @[contNetwork.scala 18:53]
    .clock(queues_50_clock),
    .reset(queues_50_reset),
    .io_addressIn_ready(queues_50_io_addressIn_ready),
    .io_addressIn_valid(queues_50_io_addressIn_valid),
    .io_addressIn_bits(queues_50_io_addressIn_bits),
    .io_addressOut_ready(queues_50_io_addressOut_ready),
    .io_addressOut_valid(queues_50_io_addressOut_valid),
    .io_addressOut_bits(queues_50_io_addressOut_bits)
  );
  contQueue queues_51 ( // @[contNetwork.scala 18:53]
    .clock(queues_51_clock),
    .reset(queues_51_reset),
    .io_addressIn_ready(queues_51_io_addressIn_ready),
    .io_addressIn_valid(queues_51_io_addressIn_valid),
    .io_addressIn_bits(queues_51_io_addressIn_bits),
    .io_addressOut_ready(queues_51_io_addressOut_ready),
    .io_addressOut_valid(queues_51_io_addressOut_valid),
    .io_addressOut_bits(queues_51_io_addressOut_bits)
  );
  contQueue queues_52 ( // @[contNetwork.scala 18:53]
    .clock(queues_52_clock),
    .reset(queues_52_reset),
    .io_addressIn_ready(queues_52_io_addressIn_ready),
    .io_addressIn_valid(queues_52_io_addressIn_valid),
    .io_addressIn_bits(queues_52_io_addressIn_bits),
    .io_addressOut_ready(queues_52_io_addressOut_ready),
    .io_addressOut_valid(queues_52_io_addressOut_valid),
    .io_addressOut_bits(queues_52_io_addressOut_bits)
  );
  contQueue queues_53 ( // @[contNetwork.scala 18:53]
    .clock(queues_53_clock),
    .reset(queues_53_reset),
    .io_addressIn_ready(queues_53_io_addressIn_ready),
    .io_addressIn_valid(queues_53_io_addressIn_valid),
    .io_addressIn_bits(queues_53_io_addressIn_bits),
    .io_addressOut_ready(queues_53_io_addressOut_ready),
    .io_addressOut_valid(queues_53_io_addressOut_valid),
    .io_addressOut_bits(queues_53_io_addressOut_bits)
  );
  contQueue queues_54 ( // @[contNetwork.scala 18:53]
    .clock(queues_54_clock),
    .reset(queues_54_reset),
    .io_addressIn_ready(queues_54_io_addressIn_ready),
    .io_addressIn_valid(queues_54_io_addressIn_valid),
    .io_addressIn_bits(queues_54_io_addressIn_bits),
    .io_addressOut_ready(queues_54_io_addressOut_ready),
    .io_addressOut_valid(queues_54_io_addressOut_valid),
    .io_addressOut_bits(queues_54_io_addressOut_bits)
  );
  contQueue queues_55 ( // @[contNetwork.scala 18:53]
    .clock(queues_55_clock),
    .reset(queues_55_reset),
    .io_addressIn_ready(queues_55_io_addressIn_ready),
    .io_addressIn_valid(queues_55_io_addressIn_valid),
    .io_addressIn_bits(queues_55_io_addressIn_bits),
    .io_addressOut_ready(queues_55_io_addressOut_ready),
    .io_addressOut_valid(queues_55_io_addressOut_valid),
    .io_addressOut_bits(queues_55_io_addressOut_bits)
  );
  contQueue queues_56 ( // @[contNetwork.scala 18:53]
    .clock(queues_56_clock),
    .reset(queues_56_reset),
    .io_addressIn_ready(queues_56_io_addressIn_ready),
    .io_addressIn_valid(queues_56_io_addressIn_valid),
    .io_addressIn_bits(queues_56_io_addressIn_bits),
    .io_addressOut_ready(queues_56_io_addressOut_ready),
    .io_addressOut_valid(queues_56_io_addressOut_valid),
    .io_addressOut_bits(queues_56_io_addressOut_bits)
  );
  contQueue queues_57 ( // @[contNetwork.scala 18:53]
    .clock(queues_57_clock),
    .reset(queues_57_reset),
    .io_addressIn_ready(queues_57_io_addressIn_ready),
    .io_addressIn_valid(queues_57_io_addressIn_valid),
    .io_addressIn_bits(queues_57_io_addressIn_bits),
    .io_addressOut_ready(queues_57_io_addressOut_ready),
    .io_addressOut_valid(queues_57_io_addressOut_valid),
    .io_addressOut_bits(queues_57_io_addressOut_bits)
  );
  contQueue queues_58 ( // @[contNetwork.scala 18:53]
    .clock(queues_58_clock),
    .reset(queues_58_reset),
    .io_addressIn_ready(queues_58_io_addressIn_ready),
    .io_addressIn_valid(queues_58_io_addressIn_valid),
    .io_addressIn_bits(queues_58_io_addressIn_bits),
    .io_addressOut_ready(queues_58_io_addressOut_ready),
    .io_addressOut_valid(queues_58_io_addressOut_valid),
    .io_addressOut_bits(queues_58_io_addressOut_bits)
  );
  contQueue queues_59 ( // @[contNetwork.scala 18:53]
    .clock(queues_59_clock),
    .reset(queues_59_reset),
    .io_addressIn_ready(queues_59_io_addressIn_ready),
    .io_addressIn_valid(queues_59_io_addressIn_valid),
    .io_addressIn_bits(queues_59_io_addressIn_bits),
    .io_addressOut_ready(queues_59_io_addressOut_ready),
    .io_addressOut_valid(queues_59_io_addressOut_valid),
    .io_addressOut_bits(queues_59_io_addressOut_bits)
  );
  contQueue queues_60 ( // @[contNetwork.scala 18:53]
    .clock(queues_60_clock),
    .reset(queues_60_reset),
    .io_addressIn_ready(queues_60_io_addressIn_ready),
    .io_addressIn_valid(queues_60_io_addressIn_valid),
    .io_addressIn_bits(queues_60_io_addressIn_bits),
    .io_addressOut_ready(queues_60_io_addressOut_ready),
    .io_addressOut_valid(queues_60_io_addressOut_valid),
    .io_addressOut_bits(queues_60_io_addressOut_bits)
  );
  contQueue queues_61 ( // @[contNetwork.scala 18:53]
    .clock(queues_61_clock),
    .reset(queues_61_reset),
    .io_addressIn_ready(queues_61_io_addressIn_ready),
    .io_addressIn_valid(queues_61_io_addressIn_valid),
    .io_addressIn_bits(queues_61_io_addressIn_bits),
    .io_addressOut_ready(queues_61_io_addressOut_ready),
    .io_addressOut_valid(queues_61_io_addressOut_valid),
    .io_addressOut_bits(queues_61_io_addressOut_bits)
  );
  contQueue queues_62 ( // @[contNetwork.scala 18:53]
    .clock(queues_62_clock),
    .reset(queues_62_reset),
    .io_addressIn_ready(queues_62_io_addressIn_ready),
    .io_addressIn_valid(queues_62_io_addressIn_valid),
    .io_addressIn_bits(queues_62_io_addressIn_bits),
    .io_addressOut_ready(queues_62_io_addressOut_ready),
    .io_addressOut_valid(queues_62_io_addressOut_valid),
    .io_addressOut_bits(queues_62_io_addressOut_bits)
  );
  contQueue queues_63 ( // @[contNetwork.scala 18:53]
    .clock(queues_63_clock),
    .reset(queues_63_reset),
    .io_addressIn_ready(queues_63_io_addressIn_ready),
    .io_addressIn_valid(queues_63_io_addressIn_valid),
    .io_addressIn_bits(queues_63_io_addressIn_bits),
    .io_addressOut_ready(queues_63_io_addressOut_ready),
    .io_addressOut_valid(queues_63_io_addressOut_valid),
    .io_addressOut_bits(queues_63_io_addressOut_bits)
  );
  assign io_connVCAS_0_ready = vcasNetworkUnits_0_io_addressIn1_ready; // @[contNetwork.scala 68:43]
  assign io_connPE_0_valid = queues_0_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_0_bits = queues_0_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_1_valid = queues_1_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_1_bits = queues_1_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_2_valid = queues_2_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_2_bits = queues_2_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_3_valid = queues_3_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_3_bits = queues_3_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_4_valid = queues_4_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_4_bits = queues_4_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_5_valid = queues_5_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_5_bits = queues_5_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_6_valid = queues_6_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_6_bits = queues_6_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_7_valid = queues_7_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_7_bits = queues_7_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_8_valid = queues_8_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_8_bits = queues_8_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_9_valid = queues_9_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_9_bits = queues_9_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_10_valid = queues_10_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_10_bits = queues_10_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_11_valid = queues_11_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_11_bits = queues_11_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_12_valid = queues_12_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_12_bits = queues_12_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_13_valid = queues_13_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_13_bits = queues_13_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_14_valid = queues_14_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_14_bits = queues_14_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_15_valid = queues_15_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_15_bits = queues_15_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_16_valid = queues_16_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_16_bits = queues_16_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_17_valid = queues_17_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_17_bits = queues_17_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_18_valid = queues_18_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_18_bits = queues_18_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_19_valid = queues_19_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_19_bits = queues_19_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_20_valid = queues_20_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_20_bits = queues_20_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_21_valid = queues_21_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_21_bits = queues_21_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_22_valid = queues_22_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_22_bits = queues_22_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_23_valid = queues_23_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_23_bits = queues_23_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_24_valid = queues_24_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_24_bits = queues_24_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_25_valid = queues_25_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_25_bits = queues_25_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_26_valid = queues_26_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_26_bits = queues_26_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_27_valid = queues_27_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_27_bits = queues_27_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_28_valid = queues_28_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_28_bits = queues_28_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_29_valid = queues_29_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_29_bits = queues_29_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_30_valid = queues_30_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_30_bits = queues_30_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_31_valid = queues_31_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_31_bits = queues_31_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_32_valid = queues_32_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_32_bits = queues_32_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_33_valid = queues_33_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_33_bits = queues_33_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_34_valid = queues_34_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_34_bits = queues_34_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_35_valid = queues_35_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_35_bits = queues_35_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_36_valid = queues_36_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_36_bits = queues_36_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_37_valid = queues_37_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_37_bits = queues_37_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_38_valid = queues_38_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_38_bits = queues_38_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_39_valid = queues_39_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_39_bits = queues_39_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_40_valid = queues_40_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_40_bits = queues_40_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_41_valid = queues_41_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_41_bits = queues_41_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_42_valid = queues_42_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_42_bits = queues_42_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_43_valid = queues_43_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_43_bits = queues_43_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_44_valid = queues_44_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_44_bits = queues_44_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_45_valid = queues_45_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_45_bits = queues_45_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_46_valid = queues_46_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_46_bits = queues_46_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_47_valid = queues_47_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_47_bits = queues_47_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_48_valid = queues_48_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_48_bits = queues_48_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_49_valid = queues_49_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_49_bits = queues_49_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_50_valid = queues_50_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_50_bits = queues_50_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_51_valid = queues_51_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_51_bits = queues_51_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_52_valid = queues_52_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_52_bits = queues_52_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_53_valid = queues_53_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_53_bits = queues_53_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_54_valid = queues_54_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_54_bits = queues_54_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_55_valid = queues_55_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_55_bits = queues_55_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_56_valid = queues_56_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_56_bits = queues_56_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_57_valid = queues_57_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_57_bits = queues_57_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_58_valid = queues_58_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_58_bits = queues_58_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_59_valid = queues_59_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_59_bits = queues_59_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_60_valid = queues_60_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_60_bits = queues_60_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_61_valid = queues_61_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_61_bits = queues_61_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_62_valid = queues_62_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_62_bits = queues_62_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign io_connPE_63_valid = queues_63_io_addressOut_valid; // @[contNetwork.scala 64:42]
  assign io_connPE_63_bits = queues_63_io_addressOut_bits; // @[contNetwork.scala 64:42]
  assign vcasNetworkUnits_0_clock = clock;
  assign vcasNetworkUnits_0_reset = reset;
  assign vcasNetworkUnits_0_io_addressIn1_valid = io_connVCAS_0_valid; // @[contNetwork.scala 68:43]
  assign vcasNetworkUnits_0_io_addressIn1_bits = io_connVCAS_0_bits; // @[contNetwork.scala 68:43]
  assign vcasNetworkUnits_0_io_addressOut_ready = networkUnits_0_io_addressIn_ready; // @[contNetwork.scala 38:67]
  assign networkUnits_0_clock = clock;
  assign networkUnits_0_reset = reset;
  assign networkUnits_0_io_addressIn_valid = vcasNetworkUnits_0_io_addressOut_valid; // @[contNetwork.scala 38:67]
  assign networkUnits_0_io_addressIn_bits = vcasNetworkUnits_0_io_addressOut_bits; // @[contNetwork.scala 38:67]
  assign networkUnits_0_io_addressOut_ready = networkUnits_1_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_0_io_casAddressOut_ready = casServers_0_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_1_clock = clock;
  assign networkUnits_1_reset = reset;
  assign networkUnits_1_io_addressIn_valid = networkUnits_0_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_1_io_addressIn_bits = networkUnits_0_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_1_io_addressOut_ready = networkUnits_2_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_1_io_casAddressOut_ready = casServers_1_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_2_clock = clock;
  assign networkUnits_2_reset = reset;
  assign networkUnits_2_io_addressIn_valid = networkUnits_1_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_2_io_addressIn_bits = networkUnits_1_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_2_io_addressOut_ready = networkUnits_3_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_2_io_casAddressOut_ready = casServers_2_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_3_clock = clock;
  assign networkUnits_3_reset = reset;
  assign networkUnits_3_io_addressIn_valid = networkUnits_2_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_3_io_addressIn_bits = networkUnits_2_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_3_io_addressOut_ready = networkUnits_4_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_3_io_casAddressOut_ready = casServers_3_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_4_clock = clock;
  assign networkUnits_4_reset = reset;
  assign networkUnits_4_io_addressIn_valid = networkUnits_3_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_4_io_addressIn_bits = networkUnits_3_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_4_io_addressOut_ready = networkUnits_5_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_4_io_casAddressOut_ready = casServers_4_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_5_clock = clock;
  assign networkUnits_5_reset = reset;
  assign networkUnits_5_io_addressIn_valid = networkUnits_4_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_5_io_addressIn_bits = networkUnits_4_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_5_io_addressOut_ready = networkUnits_6_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_5_io_casAddressOut_ready = casServers_5_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_6_clock = clock;
  assign networkUnits_6_reset = reset;
  assign networkUnits_6_io_addressIn_valid = networkUnits_5_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_6_io_addressIn_bits = networkUnits_5_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_6_io_addressOut_ready = networkUnits_7_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_6_io_casAddressOut_ready = casServers_6_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_7_clock = clock;
  assign networkUnits_7_reset = reset;
  assign networkUnits_7_io_addressIn_valid = networkUnits_6_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_7_io_addressIn_bits = networkUnits_6_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_7_io_addressOut_ready = networkUnits_8_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_7_io_casAddressOut_ready = casServers_7_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_8_clock = clock;
  assign networkUnits_8_reset = reset;
  assign networkUnits_8_io_addressIn_valid = networkUnits_7_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_8_io_addressIn_bits = networkUnits_7_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_8_io_addressOut_ready = networkUnits_9_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_8_io_casAddressOut_ready = casServers_8_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_9_clock = clock;
  assign networkUnits_9_reset = reset;
  assign networkUnits_9_io_addressIn_valid = networkUnits_8_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_9_io_addressIn_bits = networkUnits_8_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_9_io_addressOut_ready = networkUnits_10_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_9_io_casAddressOut_ready = casServers_9_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_10_clock = clock;
  assign networkUnits_10_reset = reset;
  assign networkUnits_10_io_addressIn_valid = networkUnits_9_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_10_io_addressIn_bits = networkUnits_9_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_10_io_addressOut_ready = networkUnits_11_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_10_io_casAddressOut_ready = casServers_10_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_11_clock = clock;
  assign networkUnits_11_reset = reset;
  assign networkUnits_11_io_addressIn_valid = networkUnits_10_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_11_io_addressIn_bits = networkUnits_10_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_11_io_addressOut_ready = networkUnits_12_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_11_io_casAddressOut_ready = casServers_11_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_12_clock = clock;
  assign networkUnits_12_reset = reset;
  assign networkUnits_12_io_addressIn_valid = networkUnits_11_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_12_io_addressIn_bits = networkUnits_11_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_12_io_addressOut_ready = networkUnits_13_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_12_io_casAddressOut_ready = casServers_12_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_13_clock = clock;
  assign networkUnits_13_reset = reset;
  assign networkUnits_13_io_addressIn_valid = networkUnits_12_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_13_io_addressIn_bits = networkUnits_12_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_13_io_addressOut_ready = networkUnits_14_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_13_io_casAddressOut_ready = casServers_13_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_14_clock = clock;
  assign networkUnits_14_reset = reset;
  assign networkUnits_14_io_addressIn_valid = networkUnits_13_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_14_io_addressIn_bits = networkUnits_13_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_14_io_addressOut_ready = networkUnits_15_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_14_io_casAddressOut_ready = casServers_14_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_15_clock = clock;
  assign networkUnits_15_reset = reset;
  assign networkUnits_15_io_addressIn_valid = networkUnits_14_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_15_io_addressIn_bits = networkUnits_14_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_15_io_addressOut_ready = networkUnits_16_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_15_io_casAddressOut_ready = casServers_15_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_16_clock = clock;
  assign networkUnits_16_reset = reset;
  assign networkUnits_16_io_addressIn_valid = networkUnits_15_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_16_io_addressIn_bits = networkUnits_15_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_16_io_addressOut_ready = networkUnits_17_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_16_io_casAddressOut_ready = casServers_16_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_17_clock = clock;
  assign networkUnits_17_reset = reset;
  assign networkUnits_17_io_addressIn_valid = networkUnits_16_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_17_io_addressIn_bits = networkUnits_16_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_17_io_addressOut_ready = networkUnits_18_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_17_io_casAddressOut_ready = casServers_17_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_18_clock = clock;
  assign networkUnits_18_reset = reset;
  assign networkUnits_18_io_addressIn_valid = networkUnits_17_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_18_io_addressIn_bits = networkUnits_17_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_18_io_addressOut_ready = networkUnits_19_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_18_io_casAddressOut_ready = casServers_18_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_19_clock = clock;
  assign networkUnits_19_reset = reset;
  assign networkUnits_19_io_addressIn_valid = networkUnits_18_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_19_io_addressIn_bits = networkUnits_18_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_19_io_addressOut_ready = networkUnits_20_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_19_io_casAddressOut_ready = casServers_19_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_20_clock = clock;
  assign networkUnits_20_reset = reset;
  assign networkUnits_20_io_addressIn_valid = networkUnits_19_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_20_io_addressIn_bits = networkUnits_19_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_20_io_addressOut_ready = networkUnits_21_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_20_io_casAddressOut_ready = casServers_20_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_21_clock = clock;
  assign networkUnits_21_reset = reset;
  assign networkUnits_21_io_addressIn_valid = networkUnits_20_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_21_io_addressIn_bits = networkUnits_20_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_21_io_addressOut_ready = networkUnits_22_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_21_io_casAddressOut_ready = casServers_21_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_22_clock = clock;
  assign networkUnits_22_reset = reset;
  assign networkUnits_22_io_addressIn_valid = networkUnits_21_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_22_io_addressIn_bits = networkUnits_21_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_22_io_addressOut_ready = networkUnits_23_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_22_io_casAddressOut_ready = casServers_22_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_23_clock = clock;
  assign networkUnits_23_reset = reset;
  assign networkUnits_23_io_addressIn_valid = networkUnits_22_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_23_io_addressIn_bits = networkUnits_22_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_23_io_addressOut_ready = networkUnits_24_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_23_io_casAddressOut_ready = casServers_23_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_24_clock = clock;
  assign networkUnits_24_reset = reset;
  assign networkUnits_24_io_addressIn_valid = networkUnits_23_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_24_io_addressIn_bits = networkUnits_23_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_24_io_addressOut_ready = networkUnits_25_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_24_io_casAddressOut_ready = casServers_24_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_25_clock = clock;
  assign networkUnits_25_reset = reset;
  assign networkUnits_25_io_addressIn_valid = networkUnits_24_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_25_io_addressIn_bits = networkUnits_24_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_25_io_addressOut_ready = networkUnits_26_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_25_io_casAddressOut_ready = casServers_25_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_26_clock = clock;
  assign networkUnits_26_reset = reset;
  assign networkUnits_26_io_addressIn_valid = networkUnits_25_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_26_io_addressIn_bits = networkUnits_25_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_26_io_addressOut_ready = networkUnits_27_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_26_io_casAddressOut_ready = casServers_26_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_27_clock = clock;
  assign networkUnits_27_reset = reset;
  assign networkUnits_27_io_addressIn_valid = networkUnits_26_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_27_io_addressIn_bits = networkUnits_26_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_27_io_addressOut_ready = networkUnits_28_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_27_io_casAddressOut_ready = casServers_27_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_28_clock = clock;
  assign networkUnits_28_reset = reset;
  assign networkUnits_28_io_addressIn_valid = networkUnits_27_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_28_io_addressIn_bits = networkUnits_27_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_28_io_addressOut_ready = networkUnits_29_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_28_io_casAddressOut_ready = casServers_28_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_29_clock = clock;
  assign networkUnits_29_reset = reset;
  assign networkUnits_29_io_addressIn_valid = networkUnits_28_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_29_io_addressIn_bits = networkUnits_28_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_29_io_addressOut_ready = networkUnits_30_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_29_io_casAddressOut_ready = casServers_29_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_30_clock = clock;
  assign networkUnits_30_reset = reset;
  assign networkUnits_30_io_addressIn_valid = networkUnits_29_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_30_io_addressIn_bits = networkUnits_29_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_30_io_addressOut_ready = networkUnits_31_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_30_io_casAddressOut_ready = casServers_30_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_31_clock = clock;
  assign networkUnits_31_reset = reset;
  assign networkUnits_31_io_addressIn_valid = networkUnits_30_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_31_io_addressIn_bits = networkUnits_30_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_31_io_addressOut_ready = networkUnits_32_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_31_io_casAddressOut_ready = casServers_31_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_32_clock = clock;
  assign networkUnits_32_reset = reset;
  assign networkUnits_32_io_addressIn_valid = networkUnits_31_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_32_io_addressIn_bits = networkUnits_31_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_32_io_addressOut_ready = networkUnits_33_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_32_io_casAddressOut_ready = casServers_32_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_33_clock = clock;
  assign networkUnits_33_reset = reset;
  assign networkUnits_33_io_addressIn_valid = networkUnits_32_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_33_io_addressIn_bits = networkUnits_32_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_33_io_addressOut_ready = networkUnits_34_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_33_io_casAddressOut_ready = casServers_33_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_34_clock = clock;
  assign networkUnits_34_reset = reset;
  assign networkUnits_34_io_addressIn_valid = networkUnits_33_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_34_io_addressIn_bits = networkUnits_33_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_34_io_addressOut_ready = networkUnits_35_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_34_io_casAddressOut_ready = casServers_34_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_35_clock = clock;
  assign networkUnits_35_reset = reset;
  assign networkUnits_35_io_addressIn_valid = networkUnits_34_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_35_io_addressIn_bits = networkUnits_34_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_35_io_addressOut_ready = networkUnits_36_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_35_io_casAddressOut_ready = casServers_35_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_36_clock = clock;
  assign networkUnits_36_reset = reset;
  assign networkUnits_36_io_addressIn_valid = networkUnits_35_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_36_io_addressIn_bits = networkUnits_35_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_36_io_addressOut_ready = networkUnits_37_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_36_io_casAddressOut_ready = casServers_36_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_37_clock = clock;
  assign networkUnits_37_reset = reset;
  assign networkUnits_37_io_addressIn_valid = networkUnits_36_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_37_io_addressIn_bits = networkUnits_36_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_37_io_addressOut_ready = networkUnits_38_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_37_io_casAddressOut_ready = casServers_37_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_38_clock = clock;
  assign networkUnits_38_reset = reset;
  assign networkUnits_38_io_addressIn_valid = networkUnits_37_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_38_io_addressIn_bits = networkUnits_37_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_38_io_addressOut_ready = networkUnits_39_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_38_io_casAddressOut_ready = casServers_38_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_39_clock = clock;
  assign networkUnits_39_reset = reset;
  assign networkUnits_39_io_addressIn_valid = networkUnits_38_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_39_io_addressIn_bits = networkUnits_38_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_39_io_addressOut_ready = networkUnits_40_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_39_io_casAddressOut_ready = casServers_39_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_40_clock = clock;
  assign networkUnits_40_reset = reset;
  assign networkUnits_40_io_addressIn_valid = networkUnits_39_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_40_io_addressIn_bits = networkUnits_39_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_40_io_addressOut_ready = networkUnits_41_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_40_io_casAddressOut_ready = casServers_40_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_41_clock = clock;
  assign networkUnits_41_reset = reset;
  assign networkUnits_41_io_addressIn_valid = networkUnits_40_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_41_io_addressIn_bits = networkUnits_40_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_41_io_addressOut_ready = networkUnits_42_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_41_io_casAddressOut_ready = casServers_41_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_42_clock = clock;
  assign networkUnits_42_reset = reset;
  assign networkUnits_42_io_addressIn_valid = networkUnits_41_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_42_io_addressIn_bits = networkUnits_41_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_42_io_addressOut_ready = networkUnits_43_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_42_io_casAddressOut_ready = casServers_42_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_43_clock = clock;
  assign networkUnits_43_reset = reset;
  assign networkUnits_43_io_addressIn_valid = networkUnits_42_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_43_io_addressIn_bits = networkUnits_42_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_43_io_addressOut_ready = networkUnits_44_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_43_io_casAddressOut_ready = casServers_43_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_44_clock = clock;
  assign networkUnits_44_reset = reset;
  assign networkUnits_44_io_addressIn_valid = networkUnits_43_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_44_io_addressIn_bits = networkUnits_43_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_44_io_addressOut_ready = networkUnits_45_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_44_io_casAddressOut_ready = casServers_44_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_45_clock = clock;
  assign networkUnits_45_reset = reset;
  assign networkUnits_45_io_addressIn_valid = networkUnits_44_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_45_io_addressIn_bits = networkUnits_44_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_45_io_addressOut_ready = networkUnits_46_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_45_io_casAddressOut_ready = casServers_45_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_46_clock = clock;
  assign networkUnits_46_reset = reset;
  assign networkUnits_46_io_addressIn_valid = networkUnits_45_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_46_io_addressIn_bits = networkUnits_45_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_46_io_addressOut_ready = networkUnits_47_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_46_io_casAddressOut_ready = casServers_46_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_47_clock = clock;
  assign networkUnits_47_reset = reset;
  assign networkUnits_47_io_addressIn_valid = networkUnits_46_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_47_io_addressIn_bits = networkUnits_46_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_47_io_addressOut_ready = networkUnits_48_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_47_io_casAddressOut_ready = casServers_47_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_48_clock = clock;
  assign networkUnits_48_reset = reset;
  assign networkUnits_48_io_addressIn_valid = networkUnits_47_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_48_io_addressIn_bits = networkUnits_47_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_48_io_addressOut_ready = networkUnits_49_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_48_io_casAddressOut_ready = casServers_48_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_49_clock = clock;
  assign networkUnits_49_reset = reset;
  assign networkUnits_49_io_addressIn_valid = networkUnits_48_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_49_io_addressIn_bits = networkUnits_48_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_49_io_addressOut_ready = networkUnits_50_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_49_io_casAddressOut_ready = casServers_49_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_50_clock = clock;
  assign networkUnits_50_reset = reset;
  assign networkUnits_50_io_addressIn_valid = networkUnits_49_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_50_io_addressIn_bits = networkUnits_49_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_50_io_addressOut_ready = networkUnits_51_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_50_io_casAddressOut_ready = casServers_50_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_51_clock = clock;
  assign networkUnits_51_reset = reset;
  assign networkUnits_51_io_addressIn_valid = networkUnits_50_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_51_io_addressIn_bits = networkUnits_50_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_51_io_addressOut_ready = networkUnits_52_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_51_io_casAddressOut_ready = casServers_51_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_52_clock = clock;
  assign networkUnits_52_reset = reset;
  assign networkUnits_52_io_addressIn_valid = networkUnits_51_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_52_io_addressIn_bits = networkUnits_51_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_52_io_addressOut_ready = networkUnits_53_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_52_io_casAddressOut_ready = casServers_52_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_53_clock = clock;
  assign networkUnits_53_reset = reset;
  assign networkUnits_53_io_addressIn_valid = networkUnits_52_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_53_io_addressIn_bits = networkUnits_52_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_53_io_addressOut_ready = networkUnits_54_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_53_io_casAddressOut_ready = casServers_53_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_54_clock = clock;
  assign networkUnits_54_reset = reset;
  assign networkUnits_54_io_addressIn_valid = networkUnits_53_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_54_io_addressIn_bits = networkUnits_53_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_54_io_addressOut_ready = networkUnits_55_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_54_io_casAddressOut_ready = casServers_54_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_55_clock = clock;
  assign networkUnits_55_reset = reset;
  assign networkUnits_55_io_addressIn_valid = networkUnits_54_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_55_io_addressIn_bits = networkUnits_54_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_55_io_addressOut_ready = networkUnits_56_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_55_io_casAddressOut_ready = casServers_55_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_56_clock = clock;
  assign networkUnits_56_reset = reset;
  assign networkUnits_56_io_addressIn_valid = networkUnits_55_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_56_io_addressIn_bits = networkUnits_55_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_56_io_addressOut_ready = networkUnits_57_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_56_io_casAddressOut_ready = casServers_56_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_57_clock = clock;
  assign networkUnits_57_reset = reset;
  assign networkUnits_57_io_addressIn_valid = networkUnits_56_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_57_io_addressIn_bits = networkUnits_56_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_57_io_addressOut_ready = networkUnits_58_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_57_io_casAddressOut_ready = casServers_57_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_58_clock = clock;
  assign networkUnits_58_reset = reset;
  assign networkUnits_58_io_addressIn_valid = networkUnits_57_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_58_io_addressIn_bits = networkUnits_57_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_58_io_addressOut_ready = networkUnits_59_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_58_io_casAddressOut_ready = casServers_58_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_59_clock = clock;
  assign networkUnits_59_reset = reset;
  assign networkUnits_59_io_addressIn_valid = networkUnits_58_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_59_io_addressIn_bits = networkUnits_58_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_59_io_addressOut_ready = networkUnits_60_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_59_io_casAddressOut_ready = casServers_59_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_60_clock = clock;
  assign networkUnits_60_reset = reset;
  assign networkUnits_60_io_addressIn_valid = networkUnits_59_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_60_io_addressIn_bits = networkUnits_59_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_60_io_addressOut_ready = networkUnits_61_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_60_io_casAddressOut_ready = casServers_60_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_61_clock = clock;
  assign networkUnits_61_reset = reset;
  assign networkUnits_61_io_addressIn_valid = networkUnits_60_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_61_io_addressIn_bits = networkUnits_60_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_61_io_addressOut_ready = networkUnits_62_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_61_io_casAddressOut_ready = casServers_61_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_62_clock = clock;
  assign networkUnits_62_reset = reset;
  assign networkUnits_62_io_addressIn_valid = networkUnits_61_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_62_io_addressIn_bits = networkUnits_61_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_62_io_addressOut_ready = networkUnits_63_io_addressIn_ready; // @[contNetwork.scala 50:59]
  assign networkUnits_62_io_casAddressOut_ready = casServers_62_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign networkUnits_63_clock = clock;
  assign networkUnits_63_reset = reset;
  assign networkUnits_63_io_addressIn_valid = networkUnits_62_io_addressOut_valid; // @[contNetwork.scala 50:59]
  assign networkUnits_63_io_addressIn_bits = networkUnits_62_io_addressOut_bits; // @[contNetwork.scala 50:59]
  assign networkUnits_63_io_addressOut_ready = 1'h0; // @[contNetwork.scala 57:49]
  assign networkUnits_63_io_casAddressOut_ready = casServers_63_io_addressIn_ready; // @[contNetwork.scala 62:42]
  assign casServers_0_clock = clock;
  assign casServers_0_reset = reset;
  assign casServers_0_io_addressIn_valid = networkUnits_0_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_0_io_addressIn_bits = networkUnits_0_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_0_io_addressOut_ready = queues_0_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_1_clock = clock;
  assign casServers_1_reset = reset;
  assign casServers_1_io_addressIn_valid = networkUnits_1_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_1_io_addressIn_bits = networkUnits_1_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_1_io_addressOut_ready = queues_1_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_2_clock = clock;
  assign casServers_2_reset = reset;
  assign casServers_2_io_addressIn_valid = networkUnits_2_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_2_io_addressIn_bits = networkUnits_2_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_2_io_addressOut_ready = queues_2_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_3_clock = clock;
  assign casServers_3_reset = reset;
  assign casServers_3_io_addressIn_valid = networkUnits_3_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_3_io_addressIn_bits = networkUnits_3_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_3_io_addressOut_ready = queues_3_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_4_clock = clock;
  assign casServers_4_reset = reset;
  assign casServers_4_io_addressIn_valid = networkUnits_4_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_4_io_addressIn_bits = networkUnits_4_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_4_io_addressOut_ready = queues_4_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_5_clock = clock;
  assign casServers_5_reset = reset;
  assign casServers_5_io_addressIn_valid = networkUnits_5_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_5_io_addressIn_bits = networkUnits_5_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_5_io_addressOut_ready = queues_5_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_6_clock = clock;
  assign casServers_6_reset = reset;
  assign casServers_6_io_addressIn_valid = networkUnits_6_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_6_io_addressIn_bits = networkUnits_6_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_6_io_addressOut_ready = queues_6_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_7_clock = clock;
  assign casServers_7_reset = reset;
  assign casServers_7_io_addressIn_valid = networkUnits_7_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_7_io_addressIn_bits = networkUnits_7_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_7_io_addressOut_ready = queues_7_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_8_clock = clock;
  assign casServers_8_reset = reset;
  assign casServers_8_io_addressIn_valid = networkUnits_8_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_8_io_addressIn_bits = networkUnits_8_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_8_io_addressOut_ready = queues_8_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_9_clock = clock;
  assign casServers_9_reset = reset;
  assign casServers_9_io_addressIn_valid = networkUnits_9_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_9_io_addressIn_bits = networkUnits_9_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_9_io_addressOut_ready = queues_9_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_10_clock = clock;
  assign casServers_10_reset = reset;
  assign casServers_10_io_addressIn_valid = networkUnits_10_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_10_io_addressIn_bits = networkUnits_10_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_10_io_addressOut_ready = queues_10_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_11_clock = clock;
  assign casServers_11_reset = reset;
  assign casServers_11_io_addressIn_valid = networkUnits_11_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_11_io_addressIn_bits = networkUnits_11_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_11_io_addressOut_ready = queues_11_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_12_clock = clock;
  assign casServers_12_reset = reset;
  assign casServers_12_io_addressIn_valid = networkUnits_12_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_12_io_addressIn_bits = networkUnits_12_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_12_io_addressOut_ready = queues_12_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_13_clock = clock;
  assign casServers_13_reset = reset;
  assign casServers_13_io_addressIn_valid = networkUnits_13_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_13_io_addressIn_bits = networkUnits_13_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_13_io_addressOut_ready = queues_13_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_14_clock = clock;
  assign casServers_14_reset = reset;
  assign casServers_14_io_addressIn_valid = networkUnits_14_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_14_io_addressIn_bits = networkUnits_14_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_14_io_addressOut_ready = queues_14_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_15_clock = clock;
  assign casServers_15_reset = reset;
  assign casServers_15_io_addressIn_valid = networkUnits_15_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_15_io_addressIn_bits = networkUnits_15_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_15_io_addressOut_ready = queues_15_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_16_clock = clock;
  assign casServers_16_reset = reset;
  assign casServers_16_io_addressIn_valid = networkUnits_16_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_16_io_addressIn_bits = networkUnits_16_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_16_io_addressOut_ready = queues_16_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_17_clock = clock;
  assign casServers_17_reset = reset;
  assign casServers_17_io_addressIn_valid = networkUnits_17_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_17_io_addressIn_bits = networkUnits_17_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_17_io_addressOut_ready = queues_17_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_18_clock = clock;
  assign casServers_18_reset = reset;
  assign casServers_18_io_addressIn_valid = networkUnits_18_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_18_io_addressIn_bits = networkUnits_18_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_18_io_addressOut_ready = queues_18_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_19_clock = clock;
  assign casServers_19_reset = reset;
  assign casServers_19_io_addressIn_valid = networkUnits_19_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_19_io_addressIn_bits = networkUnits_19_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_19_io_addressOut_ready = queues_19_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_20_clock = clock;
  assign casServers_20_reset = reset;
  assign casServers_20_io_addressIn_valid = networkUnits_20_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_20_io_addressIn_bits = networkUnits_20_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_20_io_addressOut_ready = queues_20_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_21_clock = clock;
  assign casServers_21_reset = reset;
  assign casServers_21_io_addressIn_valid = networkUnits_21_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_21_io_addressIn_bits = networkUnits_21_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_21_io_addressOut_ready = queues_21_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_22_clock = clock;
  assign casServers_22_reset = reset;
  assign casServers_22_io_addressIn_valid = networkUnits_22_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_22_io_addressIn_bits = networkUnits_22_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_22_io_addressOut_ready = queues_22_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_23_clock = clock;
  assign casServers_23_reset = reset;
  assign casServers_23_io_addressIn_valid = networkUnits_23_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_23_io_addressIn_bits = networkUnits_23_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_23_io_addressOut_ready = queues_23_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_24_clock = clock;
  assign casServers_24_reset = reset;
  assign casServers_24_io_addressIn_valid = networkUnits_24_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_24_io_addressIn_bits = networkUnits_24_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_24_io_addressOut_ready = queues_24_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_25_clock = clock;
  assign casServers_25_reset = reset;
  assign casServers_25_io_addressIn_valid = networkUnits_25_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_25_io_addressIn_bits = networkUnits_25_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_25_io_addressOut_ready = queues_25_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_26_clock = clock;
  assign casServers_26_reset = reset;
  assign casServers_26_io_addressIn_valid = networkUnits_26_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_26_io_addressIn_bits = networkUnits_26_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_26_io_addressOut_ready = queues_26_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_27_clock = clock;
  assign casServers_27_reset = reset;
  assign casServers_27_io_addressIn_valid = networkUnits_27_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_27_io_addressIn_bits = networkUnits_27_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_27_io_addressOut_ready = queues_27_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_28_clock = clock;
  assign casServers_28_reset = reset;
  assign casServers_28_io_addressIn_valid = networkUnits_28_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_28_io_addressIn_bits = networkUnits_28_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_28_io_addressOut_ready = queues_28_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_29_clock = clock;
  assign casServers_29_reset = reset;
  assign casServers_29_io_addressIn_valid = networkUnits_29_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_29_io_addressIn_bits = networkUnits_29_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_29_io_addressOut_ready = queues_29_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_30_clock = clock;
  assign casServers_30_reset = reset;
  assign casServers_30_io_addressIn_valid = networkUnits_30_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_30_io_addressIn_bits = networkUnits_30_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_30_io_addressOut_ready = queues_30_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_31_clock = clock;
  assign casServers_31_reset = reset;
  assign casServers_31_io_addressIn_valid = networkUnits_31_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_31_io_addressIn_bits = networkUnits_31_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_31_io_addressOut_ready = queues_31_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_32_clock = clock;
  assign casServers_32_reset = reset;
  assign casServers_32_io_addressIn_valid = networkUnits_32_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_32_io_addressIn_bits = networkUnits_32_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_32_io_addressOut_ready = queues_32_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_33_clock = clock;
  assign casServers_33_reset = reset;
  assign casServers_33_io_addressIn_valid = networkUnits_33_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_33_io_addressIn_bits = networkUnits_33_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_33_io_addressOut_ready = queues_33_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_34_clock = clock;
  assign casServers_34_reset = reset;
  assign casServers_34_io_addressIn_valid = networkUnits_34_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_34_io_addressIn_bits = networkUnits_34_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_34_io_addressOut_ready = queues_34_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_35_clock = clock;
  assign casServers_35_reset = reset;
  assign casServers_35_io_addressIn_valid = networkUnits_35_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_35_io_addressIn_bits = networkUnits_35_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_35_io_addressOut_ready = queues_35_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_36_clock = clock;
  assign casServers_36_reset = reset;
  assign casServers_36_io_addressIn_valid = networkUnits_36_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_36_io_addressIn_bits = networkUnits_36_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_36_io_addressOut_ready = queues_36_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_37_clock = clock;
  assign casServers_37_reset = reset;
  assign casServers_37_io_addressIn_valid = networkUnits_37_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_37_io_addressIn_bits = networkUnits_37_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_37_io_addressOut_ready = queues_37_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_38_clock = clock;
  assign casServers_38_reset = reset;
  assign casServers_38_io_addressIn_valid = networkUnits_38_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_38_io_addressIn_bits = networkUnits_38_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_38_io_addressOut_ready = queues_38_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_39_clock = clock;
  assign casServers_39_reset = reset;
  assign casServers_39_io_addressIn_valid = networkUnits_39_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_39_io_addressIn_bits = networkUnits_39_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_39_io_addressOut_ready = queues_39_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_40_clock = clock;
  assign casServers_40_reset = reset;
  assign casServers_40_io_addressIn_valid = networkUnits_40_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_40_io_addressIn_bits = networkUnits_40_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_40_io_addressOut_ready = queues_40_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_41_clock = clock;
  assign casServers_41_reset = reset;
  assign casServers_41_io_addressIn_valid = networkUnits_41_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_41_io_addressIn_bits = networkUnits_41_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_41_io_addressOut_ready = queues_41_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_42_clock = clock;
  assign casServers_42_reset = reset;
  assign casServers_42_io_addressIn_valid = networkUnits_42_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_42_io_addressIn_bits = networkUnits_42_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_42_io_addressOut_ready = queues_42_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_43_clock = clock;
  assign casServers_43_reset = reset;
  assign casServers_43_io_addressIn_valid = networkUnits_43_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_43_io_addressIn_bits = networkUnits_43_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_43_io_addressOut_ready = queues_43_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_44_clock = clock;
  assign casServers_44_reset = reset;
  assign casServers_44_io_addressIn_valid = networkUnits_44_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_44_io_addressIn_bits = networkUnits_44_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_44_io_addressOut_ready = queues_44_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_45_clock = clock;
  assign casServers_45_reset = reset;
  assign casServers_45_io_addressIn_valid = networkUnits_45_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_45_io_addressIn_bits = networkUnits_45_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_45_io_addressOut_ready = queues_45_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_46_clock = clock;
  assign casServers_46_reset = reset;
  assign casServers_46_io_addressIn_valid = networkUnits_46_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_46_io_addressIn_bits = networkUnits_46_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_46_io_addressOut_ready = queues_46_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_47_clock = clock;
  assign casServers_47_reset = reset;
  assign casServers_47_io_addressIn_valid = networkUnits_47_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_47_io_addressIn_bits = networkUnits_47_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_47_io_addressOut_ready = queues_47_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_48_clock = clock;
  assign casServers_48_reset = reset;
  assign casServers_48_io_addressIn_valid = networkUnits_48_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_48_io_addressIn_bits = networkUnits_48_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_48_io_addressOut_ready = queues_48_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_49_clock = clock;
  assign casServers_49_reset = reset;
  assign casServers_49_io_addressIn_valid = networkUnits_49_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_49_io_addressIn_bits = networkUnits_49_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_49_io_addressOut_ready = queues_49_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_50_clock = clock;
  assign casServers_50_reset = reset;
  assign casServers_50_io_addressIn_valid = networkUnits_50_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_50_io_addressIn_bits = networkUnits_50_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_50_io_addressOut_ready = queues_50_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_51_clock = clock;
  assign casServers_51_reset = reset;
  assign casServers_51_io_addressIn_valid = networkUnits_51_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_51_io_addressIn_bits = networkUnits_51_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_51_io_addressOut_ready = queues_51_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_52_clock = clock;
  assign casServers_52_reset = reset;
  assign casServers_52_io_addressIn_valid = networkUnits_52_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_52_io_addressIn_bits = networkUnits_52_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_52_io_addressOut_ready = queues_52_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_53_clock = clock;
  assign casServers_53_reset = reset;
  assign casServers_53_io_addressIn_valid = networkUnits_53_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_53_io_addressIn_bits = networkUnits_53_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_53_io_addressOut_ready = queues_53_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_54_clock = clock;
  assign casServers_54_reset = reset;
  assign casServers_54_io_addressIn_valid = networkUnits_54_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_54_io_addressIn_bits = networkUnits_54_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_54_io_addressOut_ready = queues_54_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_55_clock = clock;
  assign casServers_55_reset = reset;
  assign casServers_55_io_addressIn_valid = networkUnits_55_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_55_io_addressIn_bits = networkUnits_55_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_55_io_addressOut_ready = queues_55_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_56_clock = clock;
  assign casServers_56_reset = reset;
  assign casServers_56_io_addressIn_valid = networkUnits_56_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_56_io_addressIn_bits = networkUnits_56_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_56_io_addressOut_ready = queues_56_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_57_clock = clock;
  assign casServers_57_reset = reset;
  assign casServers_57_io_addressIn_valid = networkUnits_57_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_57_io_addressIn_bits = networkUnits_57_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_57_io_addressOut_ready = queues_57_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_58_clock = clock;
  assign casServers_58_reset = reset;
  assign casServers_58_io_addressIn_valid = networkUnits_58_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_58_io_addressIn_bits = networkUnits_58_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_58_io_addressOut_ready = queues_58_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_59_clock = clock;
  assign casServers_59_reset = reset;
  assign casServers_59_io_addressIn_valid = networkUnits_59_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_59_io_addressIn_bits = networkUnits_59_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_59_io_addressOut_ready = queues_59_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_60_clock = clock;
  assign casServers_60_reset = reset;
  assign casServers_60_io_addressIn_valid = networkUnits_60_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_60_io_addressIn_bits = networkUnits_60_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_60_io_addressOut_ready = queues_60_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_61_clock = clock;
  assign casServers_61_reset = reset;
  assign casServers_61_io_addressIn_valid = networkUnits_61_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_61_io_addressIn_bits = networkUnits_61_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_61_io_addressOut_ready = queues_61_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_62_clock = clock;
  assign casServers_62_reset = reset;
  assign casServers_62_io_addressIn_valid = networkUnits_62_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_62_io_addressIn_bits = networkUnits_62_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_62_io_addressOut_ready = queues_62_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign casServers_63_clock = clock;
  assign casServers_63_reset = reset;
  assign casServers_63_io_addressIn_valid = networkUnits_63_io_casAddressOut_valid; // @[contNetwork.scala 62:42]
  assign casServers_63_io_addressIn_bits = networkUnits_63_io_casAddressOut_bits; // @[contNetwork.scala 62:42]
  assign casServers_63_io_addressOut_ready = queues_63_io_addressIn_ready; // @[contNetwork.scala 63:42]
  assign queues_0_clock = clock;
  assign queues_0_reset = reset;
  assign queues_0_io_addressIn_valid = casServers_0_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_0_io_addressIn_bits = casServers_0_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_0_io_addressOut_ready = io_connPE_0_ready; // @[contNetwork.scala 64:42]
  assign queues_1_clock = clock;
  assign queues_1_reset = reset;
  assign queues_1_io_addressIn_valid = casServers_1_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_1_io_addressIn_bits = casServers_1_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_1_io_addressOut_ready = io_connPE_1_ready; // @[contNetwork.scala 64:42]
  assign queues_2_clock = clock;
  assign queues_2_reset = reset;
  assign queues_2_io_addressIn_valid = casServers_2_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_2_io_addressIn_bits = casServers_2_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_2_io_addressOut_ready = io_connPE_2_ready; // @[contNetwork.scala 64:42]
  assign queues_3_clock = clock;
  assign queues_3_reset = reset;
  assign queues_3_io_addressIn_valid = casServers_3_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_3_io_addressIn_bits = casServers_3_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_3_io_addressOut_ready = io_connPE_3_ready; // @[contNetwork.scala 64:42]
  assign queues_4_clock = clock;
  assign queues_4_reset = reset;
  assign queues_4_io_addressIn_valid = casServers_4_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_4_io_addressIn_bits = casServers_4_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_4_io_addressOut_ready = io_connPE_4_ready; // @[contNetwork.scala 64:42]
  assign queues_5_clock = clock;
  assign queues_5_reset = reset;
  assign queues_5_io_addressIn_valid = casServers_5_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_5_io_addressIn_bits = casServers_5_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_5_io_addressOut_ready = io_connPE_5_ready; // @[contNetwork.scala 64:42]
  assign queues_6_clock = clock;
  assign queues_6_reset = reset;
  assign queues_6_io_addressIn_valid = casServers_6_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_6_io_addressIn_bits = casServers_6_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_6_io_addressOut_ready = io_connPE_6_ready; // @[contNetwork.scala 64:42]
  assign queues_7_clock = clock;
  assign queues_7_reset = reset;
  assign queues_7_io_addressIn_valid = casServers_7_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_7_io_addressIn_bits = casServers_7_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_7_io_addressOut_ready = io_connPE_7_ready; // @[contNetwork.scala 64:42]
  assign queues_8_clock = clock;
  assign queues_8_reset = reset;
  assign queues_8_io_addressIn_valid = casServers_8_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_8_io_addressIn_bits = casServers_8_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_8_io_addressOut_ready = io_connPE_8_ready; // @[contNetwork.scala 64:42]
  assign queues_9_clock = clock;
  assign queues_9_reset = reset;
  assign queues_9_io_addressIn_valid = casServers_9_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_9_io_addressIn_bits = casServers_9_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_9_io_addressOut_ready = io_connPE_9_ready; // @[contNetwork.scala 64:42]
  assign queues_10_clock = clock;
  assign queues_10_reset = reset;
  assign queues_10_io_addressIn_valid = casServers_10_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_10_io_addressIn_bits = casServers_10_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_10_io_addressOut_ready = io_connPE_10_ready; // @[contNetwork.scala 64:42]
  assign queues_11_clock = clock;
  assign queues_11_reset = reset;
  assign queues_11_io_addressIn_valid = casServers_11_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_11_io_addressIn_bits = casServers_11_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_11_io_addressOut_ready = io_connPE_11_ready; // @[contNetwork.scala 64:42]
  assign queues_12_clock = clock;
  assign queues_12_reset = reset;
  assign queues_12_io_addressIn_valid = casServers_12_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_12_io_addressIn_bits = casServers_12_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_12_io_addressOut_ready = io_connPE_12_ready; // @[contNetwork.scala 64:42]
  assign queues_13_clock = clock;
  assign queues_13_reset = reset;
  assign queues_13_io_addressIn_valid = casServers_13_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_13_io_addressIn_bits = casServers_13_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_13_io_addressOut_ready = io_connPE_13_ready; // @[contNetwork.scala 64:42]
  assign queues_14_clock = clock;
  assign queues_14_reset = reset;
  assign queues_14_io_addressIn_valid = casServers_14_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_14_io_addressIn_bits = casServers_14_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_14_io_addressOut_ready = io_connPE_14_ready; // @[contNetwork.scala 64:42]
  assign queues_15_clock = clock;
  assign queues_15_reset = reset;
  assign queues_15_io_addressIn_valid = casServers_15_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_15_io_addressIn_bits = casServers_15_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_15_io_addressOut_ready = io_connPE_15_ready; // @[contNetwork.scala 64:42]
  assign queues_16_clock = clock;
  assign queues_16_reset = reset;
  assign queues_16_io_addressIn_valid = casServers_16_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_16_io_addressIn_bits = casServers_16_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_16_io_addressOut_ready = io_connPE_16_ready; // @[contNetwork.scala 64:42]
  assign queues_17_clock = clock;
  assign queues_17_reset = reset;
  assign queues_17_io_addressIn_valid = casServers_17_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_17_io_addressIn_bits = casServers_17_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_17_io_addressOut_ready = io_connPE_17_ready; // @[contNetwork.scala 64:42]
  assign queues_18_clock = clock;
  assign queues_18_reset = reset;
  assign queues_18_io_addressIn_valid = casServers_18_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_18_io_addressIn_bits = casServers_18_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_18_io_addressOut_ready = io_connPE_18_ready; // @[contNetwork.scala 64:42]
  assign queues_19_clock = clock;
  assign queues_19_reset = reset;
  assign queues_19_io_addressIn_valid = casServers_19_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_19_io_addressIn_bits = casServers_19_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_19_io_addressOut_ready = io_connPE_19_ready; // @[contNetwork.scala 64:42]
  assign queues_20_clock = clock;
  assign queues_20_reset = reset;
  assign queues_20_io_addressIn_valid = casServers_20_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_20_io_addressIn_bits = casServers_20_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_20_io_addressOut_ready = io_connPE_20_ready; // @[contNetwork.scala 64:42]
  assign queues_21_clock = clock;
  assign queues_21_reset = reset;
  assign queues_21_io_addressIn_valid = casServers_21_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_21_io_addressIn_bits = casServers_21_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_21_io_addressOut_ready = io_connPE_21_ready; // @[contNetwork.scala 64:42]
  assign queues_22_clock = clock;
  assign queues_22_reset = reset;
  assign queues_22_io_addressIn_valid = casServers_22_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_22_io_addressIn_bits = casServers_22_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_22_io_addressOut_ready = io_connPE_22_ready; // @[contNetwork.scala 64:42]
  assign queues_23_clock = clock;
  assign queues_23_reset = reset;
  assign queues_23_io_addressIn_valid = casServers_23_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_23_io_addressIn_bits = casServers_23_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_23_io_addressOut_ready = io_connPE_23_ready; // @[contNetwork.scala 64:42]
  assign queues_24_clock = clock;
  assign queues_24_reset = reset;
  assign queues_24_io_addressIn_valid = casServers_24_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_24_io_addressIn_bits = casServers_24_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_24_io_addressOut_ready = io_connPE_24_ready; // @[contNetwork.scala 64:42]
  assign queues_25_clock = clock;
  assign queues_25_reset = reset;
  assign queues_25_io_addressIn_valid = casServers_25_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_25_io_addressIn_bits = casServers_25_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_25_io_addressOut_ready = io_connPE_25_ready; // @[contNetwork.scala 64:42]
  assign queues_26_clock = clock;
  assign queues_26_reset = reset;
  assign queues_26_io_addressIn_valid = casServers_26_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_26_io_addressIn_bits = casServers_26_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_26_io_addressOut_ready = io_connPE_26_ready; // @[contNetwork.scala 64:42]
  assign queues_27_clock = clock;
  assign queues_27_reset = reset;
  assign queues_27_io_addressIn_valid = casServers_27_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_27_io_addressIn_bits = casServers_27_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_27_io_addressOut_ready = io_connPE_27_ready; // @[contNetwork.scala 64:42]
  assign queues_28_clock = clock;
  assign queues_28_reset = reset;
  assign queues_28_io_addressIn_valid = casServers_28_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_28_io_addressIn_bits = casServers_28_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_28_io_addressOut_ready = io_connPE_28_ready; // @[contNetwork.scala 64:42]
  assign queues_29_clock = clock;
  assign queues_29_reset = reset;
  assign queues_29_io_addressIn_valid = casServers_29_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_29_io_addressIn_bits = casServers_29_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_29_io_addressOut_ready = io_connPE_29_ready; // @[contNetwork.scala 64:42]
  assign queues_30_clock = clock;
  assign queues_30_reset = reset;
  assign queues_30_io_addressIn_valid = casServers_30_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_30_io_addressIn_bits = casServers_30_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_30_io_addressOut_ready = io_connPE_30_ready; // @[contNetwork.scala 64:42]
  assign queues_31_clock = clock;
  assign queues_31_reset = reset;
  assign queues_31_io_addressIn_valid = casServers_31_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_31_io_addressIn_bits = casServers_31_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_31_io_addressOut_ready = io_connPE_31_ready; // @[contNetwork.scala 64:42]
  assign queues_32_clock = clock;
  assign queues_32_reset = reset;
  assign queues_32_io_addressIn_valid = casServers_32_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_32_io_addressIn_bits = casServers_32_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_32_io_addressOut_ready = io_connPE_32_ready; // @[contNetwork.scala 64:42]
  assign queues_33_clock = clock;
  assign queues_33_reset = reset;
  assign queues_33_io_addressIn_valid = casServers_33_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_33_io_addressIn_bits = casServers_33_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_33_io_addressOut_ready = io_connPE_33_ready; // @[contNetwork.scala 64:42]
  assign queues_34_clock = clock;
  assign queues_34_reset = reset;
  assign queues_34_io_addressIn_valid = casServers_34_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_34_io_addressIn_bits = casServers_34_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_34_io_addressOut_ready = io_connPE_34_ready; // @[contNetwork.scala 64:42]
  assign queues_35_clock = clock;
  assign queues_35_reset = reset;
  assign queues_35_io_addressIn_valid = casServers_35_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_35_io_addressIn_bits = casServers_35_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_35_io_addressOut_ready = io_connPE_35_ready; // @[contNetwork.scala 64:42]
  assign queues_36_clock = clock;
  assign queues_36_reset = reset;
  assign queues_36_io_addressIn_valid = casServers_36_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_36_io_addressIn_bits = casServers_36_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_36_io_addressOut_ready = io_connPE_36_ready; // @[contNetwork.scala 64:42]
  assign queues_37_clock = clock;
  assign queues_37_reset = reset;
  assign queues_37_io_addressIn_valid = casServers_37_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_37_io_addressIn_bits = casServers_37_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_37_io_addressOut_ready = io_connPE_37_ready; // @[contNetwork.scala 64:42]
  assign queues_38_clock = clock;
  assign queues_38_reset = reset;
  assign queues_38_io_addressIn_valid = casServers_38_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_38_io_addressIn_bits = casServers_38_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_38_io_addressOut_ready = io_connPE_38_ready; // @[contNetwork.scala 64:42]
  assign queues_39_clock = clock;
  assign queues_39_reset = reset;
  assign queues_39_io_addressIn_valid = casServers_39_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_39_io_addressIn_bits = casServers_39_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_39_io_addressOut_ready = io_connPE_39_ready; // @[contNetwork.scala 64:42]
  assign queues_40_clock = clock;
  assign queues_40_reset = reset;
  assign queues_40_io_addressIn_valid = casServers_40_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_40_io_addressIn_bits = casServers_40_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_40_io_addressOut_ready = io_connPE_40_ready; // @[contNetwork.scala 64:42]
  assign queues_41_clock = clock;
  assign queues_41_reset = reset;
  assign queues_41_io_addressIn_valid = casServers_41_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_41_io_addressIn_bits = casServers_41_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_41_io_addressOut_ready = io_connPE_41_ready; // @[contNetwork.scala 64:42]
  assign queues_42_clock = clock;
  assign queues_42_reset = reset;
  assign queues_42_io_addressIn_valid = casServers_42_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_42_io_addressIn_bits = casServers_42_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_42_io_addressOut_ready = io_connPE_42_ready; // @[contNetwork.scala 64:42]
  assign queues_43_clock = clock;
  assign queues_43_reset = reset;
  assign queues_43_io_addressIn_valid = casServers_43_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_43_io_addressIn_bits = casServers_43_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_43_io_addressOut_ready = io_connPE_43_ready; // @[contNetwork.scala 64:42]
  assign queues_44_clock = clock;
  assign queues_44_reset = reset;
  assign queues_44_io_addressIn_valid = casServers_44_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_44_io_addressIn_bits = casServers_44_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_44_io_addressOut_ready = io_connPE_44_ready; // @[contNetwork.scala 64:42]
  assign queues_45_clock = clock;
  assign queues_45_reset = reset;
  assign queues_45_io_addressIn_valid = casServers_45_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_45_io_addressIn_bits = casServers_45_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_45_io_addressOut_ready = io_connPE_45_ready; // @[contNetwork.scala 64:42]
  assign queues_46_clock = clock;
  assign queues_46_reset = reset;
  assign queues_46_io_addressIn_valid = casServers_46_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_46_io_addressIn_bits = casServers_46_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_46_io_addressOut_ready = io_connPE_46_ready; // @[contNetwork.scala 64:42]
  assign queues_47_clock = clock;
  assign queues_47_reset = reset;
  assign queues_47_io_addressIn_valid = casServers_47_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_47_io_addressIn_bits = casServers_47_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_47_io_addressOut_ready = io_connPE_47_ready; // @[contNetwork.scala 64:42]
  assign queues_48_clock = clock;
  assign queues_48_reset = reset;
  assign queues_48_io_addressIn_valid = casServers_48_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_48_io_addressIn_bits = casServers_48_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_48_io_addressOut_ready = io_connPE_48_ready; // @[contNetwork.scala 64:42]
  assign queues_49_clock = clock;
  assign queues_49_reset = reset;
  assign queues_49_io_addressIn_valid = casServers_49_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_49_io_addressIn_bits = casServers_49_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_49_io_addressOut_ready = io_connPE_49_ready; // @[contNetwork.scala 64:42]
  assign queues_50_clock = clock;
  assign queues_50_reset = reset;
  assign queues_50_io_addressIn_valid = casServers_50_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_50_io_addressIn_bits = casServers_50_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_50_io_addressOut_ready = io_connPE_50_ready; // @[contNetwork.scala 64:42]
  assign queues_51_clock = clock;
  assign queues_51_reset = reset;
  assign queues_51_io_addressIn_valid = casServers_51_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_51_io_addressIn_bits = casServers_51_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_51_io_addressOut_ready = io_connPE_51_ready; // @[contNetwork.scala 64:42]
  assign queues_52_clock = clock;
  assign queues_52_reset = reset;
  assign queues_52_io_addressIn_valid = casServers_52_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_52_io_addressIn_bits = casServers_52_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_52_io_addressOut_ready = io_connPE_52_ready; // @[contNetwork.scala 64:42]
  assign queues_53_clock = clock;
  assign queues_53_reset = reset;
  assign queues_53_io_addressIn_valid = casServers_53_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_53_io_addressIn_bits = casServers_53_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_53_io_addressOut_ready = io_connPE_53_ready; // @[contNetwork.scala 64:42]
  assign queues_54_clock = clock;
  assign queues_54_reset = reset;
  assign queues_54_io_addressIn_valid = casServers_54_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_54_io_addressIn_bits = casServers_54_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_54_io_addressOut_ready = io_connPE_54_ready; // @[contNetwork.scala 64:42]
  assign queues_55_clock = clock;
  assign queues_55_reset = reset;
  assign queues_55_io_addressIn_valid = casServers_55_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_55_io_addressIn_bits = casServers_55_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_55_io_addressOut_ready = io_connPE_55_ready; // @[contNetwork.scala 64:42]
  assign queues_56_clock = clock;
  assign queues_56_reset = reset;
  assign queues_56_io_addressIn_valid = casServers_56_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_56_io_addressIn_bits = casServers_56_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_56_io_addressOut_ready = io_connPE_56_ready; // @[contNetwork.scala 64:42]
  assign queues_57_clock = clock;
  assign queues_57_reset = reset;
  assign queues_57_io_addressIn_valid = casServers_57_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_57_io_addressIn_bits = casServers_57_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_57_io_addressOut_ready = io_connPE_57_ready; // @[contNetwork.scala 64:42]
  assign queues_58_clock = clock;
  assign queues_58_reset = reset;
  assign queues_58_io_addressIn_valid = casServers_58_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_58_io_addressIn_bits = casServers_58_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_58_io_addressOut_ready = io_connPE_58_ready; // @[contNetwork.scala 64:42]
  assign queues_59_clock = clock;
  assign queues_59_reset = reset;
  assign queues_59_io_addressIn_valid = casServers_59_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_59_io_addressIn_bits = casServers_59_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_59_io_addressOut_ready = io_connPE_59_ready; // @[contNetwork.scala 64:42]
  assign queues_60_clock = clock;
  assign queues_60_reset = reset;
  assign queues_60_io_addressIn_valid = casServers_60_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_60_io_addressIn_bits = casServers_60_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_60_io_addressOut_ready = io_connPE_60_ready; // @[contNetwork.scala 64:42]
  assign queues_61_clock = clock;
  assign queues_61_reset = reset;
  assign queues_61_io_addressIn_valid = casServers_61_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_61_io_addressIn_bits = casServers_61_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_61_io_addressOut_ready = io_connPE_61_ready; // @[contNetwork.scala 64:42]
  assign queues_62_clock = clock;
  assign queues_62_reset = reset;
  assign queues_62_io_addressIn_valid = casServers_62_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_62_io_addressIn_bits = casServers_62_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_62_io_addressOut_ready = io_connPE_62_ready; // @[contNetwork.scala 64:42]
  assign queues_63_clock = clock;
  assign queues_63_reset = reset;
  assign queues_63_io_addressIn_valid = casServers_63_io_addressOut_valid; // @[contNetwork.scala 63:42]
  assign queues_63_io_addressIn_bits = casServers_63_io_addressOut_bits; // @[contNetwork.scala 63:42]
  assign queues_63_io_addressOut_ready = io_connPE_63_ready; // @[contNetwork.scala 64:42]
endmodule
module virtContAddrServer(
  input         clock,
  input         reset,
  input         io_dataOut_ready,
  output        io_dataOut_valid,
  output [63:0] io_dataOut_bits,
  output        io_axi_mgmt_ARREADY,
  input         io_axi_mgmt_ARVALID,
  input  [5:0]  io_axi_mgmt_ARADDR,
  input         io_axi_mgmt_RREADY,
  output        io_axi_mgmt_RVALID,
  output [63:0] io_axi_mgmt_RDATA,
  output        io_axi_mgmt_AWREADY,
  input         io_axi_mgmt_AWVALID,
  input  [5:0]  io_axi_mgmt_AWADDR,
  output        io_axi_mgmt_WREADY,
  input         io_axi_mgmt_WVALID,
  input  [63:0] io_axi_mgmt_WDATA,
  input  [7:0]  io_axi_mgmt_WSTRB,
  input         io_axi_mgmt_BREADY,
  output        io_axi_mgmt_BVALID,
  input         io_read_address_ready,
  output        io_read_address_valid,
  output [63:0] io_read_address_bits,
  output        io_read_data_ready,
  input         io_read_data_valid,
  input  [63:0] io_read_data_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire  rdReq__deq_clock; // @[Decoupled.scala 377:21]
  wire  rdReq__deq_reset; // @[Decoupled.scala 377:21]
  wire  rdReq__deq_io_enq_ready; // @[Decoupled.scala 377:21]
  wire  rdReq__deq_io_enq_valid; // @[Decoupled.scala 377:21]
  wire [5:0] rdReq__deq_io_enq_bits_addr; // @[Decoupled.scala 377:21]
  wire  rdReq__deq_io_deq_ready; // @[Decoupled.scala 377:21]
  wire  rdReq__deq_io_deq_valid; // @[Decoupled.scala 377:21]
  wire [5:0] rdReq__deq_io_deq_bits_addr; // @[Decoupled.scala 377:21]
  wire  wrReq__deq_clock; // @[Decoupled.scala 377:21]
  wire  wrReq__deq_reset; // @[Decoupled.scala 377:21]
  wire  wrReq__deq_io_enq_ready; // @[Decoupled.scala 377:21]
  wire  wrReq__deq_io_enq_valid; // @[Decoupled.scala 377:21]
  wire [5:0] wrReq__deq_io_enq_bits_addr; // @[Decoupled.scala 377:21]
  wire  wrReq__deq_io_deq_ready; // @[Decoupled.scala 377:21]
  wire  wrReq__deq_io_deq_valid; // @[Decoupled.scala 377:21]
  wire [5:0] wrReq__deq_io_deq_bits_addr; // @[Decoupled.scala 377:21]
  wire  wrReqData__deq_clock; // @[Decoupled.scala 377:21]
  wire  wrReqData__deq_reset; // @[Decoupled.scala 377:21]
  wire  wrReqData__deq_io_enq_ready; // @[Decoupled.scala 377:21]
  wire  wrReqData__deq_io_enq_valid; // @[Decoupled.scala 377:21]
  wire [63:0] wrReqData__deq_io_enq_bits_data; // @[Decoupled.scala 377:21]
  wire [7:0] wrReqData__deq_io_enq_bits_strb; // @[Decoupled.scala 377:21]
  wire  wrReqData__deq_io_deq_ready; // @[Decoupled.scala 377:21]
  wire  wrReqData__deq_io_deq_valid; // @[Decoupled.scala 377:21]
  wire [63:0] wrReqData__deq_io_deq_bits_data; // @[Decoupled.scala 377:21]
  wire [7:0] wrReqData__deq_io_deq_bits_strb; // @[Decoupled.scala 377:21]
  wire  rdReq__valid = rdReq__deq_io_deq_valid; // @[Decoupled.scala 417:19 419:15]
  wire  rdReq = rdReq__valid & io_axi_mgmt_RREADY; // @[RegisterBlock.scala 210:44]
  wire [5:0] rdReq__bits_addr = rdReq__deq_io_deq_bits_addr; // @[Decoupled.scala 417:19 418:14]
  wire [5:0] rdAddr = rdReq__bits_addr & 6'h38; // @[RegisterBlock.scala 214:48]
  wire  wrReq__valid = wrReq__deq_io_deq_valid; // @[Decoupled.scala 417:19 419:15]
  wire  wrReqData__valid = wrReqData__deq_io_deq_valid; // @[Decoupled.scala 417:19 419:15]
  wire  wrReq = wrReq__valid & wrReqData__valid & io_axi_mgmt_BREADY; // @[RegisterBlock.scala 241:63]
  wire [5:0] wrReq__bits_addr = wrReq__deq_io_deq_bits_addr; // @[Decoupled.scala 417:19 418:14]
  wire [5:0] wrAddr = wrReq__bits_addr & 6'h38; // @[RegisterBlock.scala 243:48]
  reg [63:0] rAddr; // @[virtContAddrServer.scala 37:49]
  reg [63:0] rPause; // @[virtContAddrServer.scala 38:49]
  reg [63:0] avaialbleSize; // @[virtContAddrServer.scala 39:49]
  reg [2:0] stateReg; // @[virtContAddrServer.scala 40:49]
  wire [63:0] index = avaialbleSize - 64'h10; // @[virtContAddrServer.scala 42:56]
  reg [63:0] continuationsRegisters_0; // @[virtContAddrServer.scala 43:49]
  reg [63:0] continuationsRegisters_1; // @[virtContAddrServer.scala 43:49]
  reg [63:0] continuationsRegisters_2; // @[virtContAddrServer.scala 43:49]
  reg [63:0] continuationsRegisters_3; // @[virtContAddrServer.scala 43:49]
  reg [63:0] continuationsRegisters_4; // @[virtContAddrServer.scala 43:49]
  reg [63:0] continuationsRegisters_5; // @[virtContAddrServer.scala 43:49]
  reg [63:0] continuationsRegisters_6; // @[virtContAddrServer.scala 43:49]
  reg [63:0] continuationsRegisters_7; // @[virtContAddrServer.scala 43:49]
  reg [63:0] continuationsRegisters_8; // @[virtContAddrServer.scala 43:49]
  reg [63:0] continuationsRegisters_9; // @[virtContAddrServer.scala 43:49]
  reg [63:0] continuationsRegisters_10; // @[virtContAddrServer.scala 43:49]
  reg [63:0] continuationsRegisters_11; // @[virtContAddrServer.scala 43:49]
  reg [63:0] continuationsRegisters_12; // @[virtContAddrServer.scala 43:49]
  reg [63:0] continuationsRegisters_13; // @[virtContAddrServer.scala 43:49]
  reg [63:0] continuationsRegisters_14; // @[virtContAddrServer.scala 43:49]
  reg [63:0] continuationsRegisters_15; // @[virtContAddrServer.scala 43:49]
  reg [3:0] burstCounter; // @[virtContAddrServer.scala 44:49]
  wire [63:0] _GEN_1 = avaialbleSize >= 64'h10 ? rPause : 64'hffffffffffffffff; // @[virtContAddrServer.scala 38:49 52:52 56:22]
  wire  _T_2 = stateReg == 3'h1; // @[virtContAddrServer.scala 58:25]
  wire  _T_3 = stateReg == 3'h2; // @[virtContAddrServer.scala 63:25]
  wire [63:0] _GEN_4 = 4'h0 == burstCounter ? io_read_data_bits : continuationsRegisters_0; // @[virtContAddrServer.scala 43:49 65:{50,50}]
  wire [63:0] _GEN_5 = 4'h1 == burstCounter ? io_read_data_bits : continuationsRegisters_1; // @[virtContAddrServer.scala 43:49 65:{50,50}]
  wire [63:0] _GEN_6 = 4'h2 == burstCounter ? io_read_data_bits : continuationsRegisters_2; // @[virtContAddrServer.scala 43:49 65:{50,50}]
  wire [63:0] _GEN_7 = 4'h3 == burstCounter ? io_read_data_bits : continuationsRegisters_3; // @[virtContAddrServer.scala 43:49 65:{50,50}]
  wire [63:0] _GEN_8 = 4'h4 == burstCounter ? io_read_data_bits : continuationsRegisters_4; // @[virtContAddrServer.scala 43:49 65:{50,50}]
  wire [63:0] _GEN_9 = 4'h5 == burstCounter ? io_read_data_bits : continuationsRegisters_5; // @[virtContAddrServer.scala 43:49 65:{50,50}]
  wire [63:0] _GEN_10 = 4'h6 == burstCounter ? io_read_data_bits : continuationsRegisters_6; // @[virtContAddrServer.scala 43:49 65:{50,50}]
  wire [63:0] _GEN_11 = 4'h7 == burstCounter ? io_read_data_bits : continuationsRegisters_7; // @[virtContAddrServer.scala 43:49 65:{50,50}]
  wire [63:0] _GEN_12 = 4'h8 == burstCounter ? io_read_data_bits : continuationsRegisters_8; // @[virtContAddrServer.scala 43:49 65:{50,50}]
  wire [63:0] _GEN_13 = 4'h9 == burstCounter ? io_read_data_bits : continuationsRegisters_9; // @[virtContAddrServer.scala 43:49 65:{50,50}]
  wire [63:0] _GEN_14 = 4'ha == burstCounter ? io_read_data_bits : continuationsRegisters_10; // @[virtContAddrServer.scala 43:49 65:{50,50}]
  wire [63:0] _GEN_15 = 4'hb == burstCounter ? io_read_data_bits : continuationsRegisters_11; // @[virtContAddrServer.scala 43:49 65:{50,50}]
  wire [63:0] _GEN_16 = 4'hc == burstCounter ? io_read_data_bits : continuationsRegisters_12; // @[virtContAddrServer.scala 43:49 65:{50,50}]
  wire [63:0] _GEN_17 = 4'hd == burstCounter ? io_read_data_bits : continuationsRegisters_13; // @[virtContAddrServer.scala 43:49 65:{50,50}]
  wire [63:0] _GEN_18 = 4'he == burstCounter ? io_read_data_bits : continuationsRegisters_14; // @[virtContAddrServer.scala 43:49 65:{50,50}]
  wire [63:0] _GEN_19 = 4'hf == burstCounter ? io_read_data_bits : continuationsRegisters_15; // @[virtContAddrServer.scala 43:49 65:{50,50}]
  wire [3:0] _burstCounter_T_1 = burstCounter - 4'h1; // @[virtContAddrServer.scala 66:66]
  wire [63:0] _avaialbleSize_T_1 = avaialbleSize - 64'h1; // @[virtContAddrServer.scala 67:44]
  wire [63:0] _GEN_20 = io_read_data_valid ? _GEN_4 : continuationsRegisters_0; // @[virtContAddrServer.scala 64:33 43:49]
  wire [63:0] _GEN_21 = io_read_data_valid ? _GEN_5 : continuationsRegisters_1; // @[virtContAddrServer.scala 64:33 43:49]
  wire [63:0] _GEN_22 = io_read_data_valid ? _GEN_6 : continuationsRegisters_2; // @[virtContAddrServer.scala 64:33 43:49]
  wire [63:0] _GEN_23 = io_read_data_valid ? _GEN_7 : continuationsRegisters_3; // @[virtContAddrServer.scala 64:33 43:49]
  wire [63:0] _GEN_24 = io_read_data_valid ? _GEN_8 : continuationsRegisters_4; // @[virtContAddrServer.scala 64:33 43:49]
  wire [63:0] _GEN_25 = io_read_data_valid ? _GEN_9 : continuationsRegisters_5; // @[virtContAddrServer.scala 64:33 43:49]
  wire [63:0] _GEN_26 = io_read_data_valid ? _GEN_10 : continuationsRegisters_6; // @[virtContAddrServer.scala 64:33 43:49]
  wire [63:0] _GEN_27 = io_read_data_valid ? _GEN_11 : continuationsRegisters_7; // @[virtContAddrServer.scala 64:33 43:49]
  wire [63:0] _GEN_28 = io_read_data_valid ? _GEN_12 : continuationsRegisters_8; // @[virtContAddrServer.scala 64:33 43:49]
  wire [63:0] _GEN_29 = io_read_data_valid ? _GEN_13 : continuationsRegisters_9; // @[virtContAddrServer.scala 64:33 43:49]
  wire [63:0] _GEN_30 = io_read_data_valid ? _GEN_14 : continuationsRegisters_10; // @[virtContAddrServer.scala 64:33 43:49]
  wire [63:0] _GEN_31 = io_read_data_valid ? _GEN_15 : continuationsRegisters_11; // @[virtContAddrServer.scala 64:33 43:49]
  wire [63:0] _GEN_32 = io_read_data_valid ? _GEN_16 : continuationsRegisters_12; // @[virtContAddrServer.scala 64:33 43:49]
  wire [63:0] _GEN_33 = io_read_data_valid ? _GEN_17 : continuationsRegisters_13; // @[virtContAddrServer.scala 64:33 43:49]
  wire [63:0] _GEN_34 = io_read_data_valid ? _GEN_18 : continuationsRegisters_14; // @[virtContAddrServer.scala 64:33 43:49]
  wire [63:0] _GEN_35 = io_read_data_valid ? _GEN_19 : continuationsRegisters_15; // @[virtContAddrServer.scala 64:33 43:49]
  wire [3:0] _GEN_36 = io_read_data_valid ? _burstCounter_T_1 : burstCounter; // @[virtContAddrServer.scala 64:33 44:49 66:50]
  wire [63:0] _GEN_37 = io_read_data_valid ? _avaialbleSize_T_1 : avaialbleSize; // @[virtContAddrServer.scala 64:33 67:27 39:49]
  wire  _T_4 = burstCounter == 4'h0; // @[virtContAddrServer.scala 70:27]
  wire [2:0] _GEN_38 = burstCounter == 4'h0 & io_read_data_valid ? 3'h3 : stateReg; // @[virtContAddrServer.scala 70:57 71:27 40:49]
  wire [63:0] _GEN_39 = burstCounter == 4'h0 & io_read_data_valid ? index : _GEN_37; // @[virtContAddrServer.scala 70:57 72:27]
  wire [3:0] _GEN_40 = burstCounter == 4'h0 & io_read_data_valid ? 4'hf : _GEN_36; // @[virtContAddrServer.scala 70:57 73:27]
  wire  _T_6 = stateReg == 3'h3; // @[virtContAddrServer.scala 76:25]
  wire [3:0] _GEN_41 = io_dataOut_ready ? _burstCounter_T_1 : burstCounter; // @[virtContAddrServer.scala 77:31 78:26 44:49]
  wire [2:0] _GEN_42 = _T_4 & io_dataOut_ready ? 3'h0 : stateReg; // @[virtContAddrServer.scala 80:55 81:22 40:49]
  wire [2:0] _GEN_43 = rPause == 64'h0 ? 3'h0 : stateReg; // @[virtContAddrServer.scala 85:33 86:22 40:49]
  wire [2:0] _GEN_44 = stateReg == 3'h4 ? _GEN_43 : stateReg; // @[virtContAddrServer.scala 84:46 40:49]
  wire [3:0] _GEN_45 = stateReg == 3'h3 ? _GEN_41 : burstCounter; // @[virtContAddrServer.scala 76:44 44:49]
  wire [2:0] _GEN_46 = stateReg == 3'h3 ? _GEN_42 : _GEN_44; // @[virtContAddrServer.scala 76:44]
  wire [63:0] _GEN_64 = stateReg == 3'h2 ? _GEN_39 : avaialbleSize; // @[virtContAddrServer.scala 63:44 39:49]
  wire [63:0] _GEN_84 = stateReg == 3'h1 ? avaialbleSize : _GEN_64; // @[virtContAddrServer.scala 39:49 58:54]
  wire [63:0] _GEN_86 = stateReg == 3'h0 ? _GEN_1 : rPause; // @[virtContAddrServer.scala 51:34 38:49]
  wire [63:0] _GEN_104 = stateReg == 3'h0 ? avaialbleSize : _GEN_84; // @[virtContAddrServer.scala 51:34 39:49]
  wire  _GEN_107 = _T_3 ? 1'h0 : _T_6; // @[virtContAddrServer.scala 92:27 98:44]
  wire [66:0] _io_read_address_bits_T = {index, 3'h0}; // @[virtContAddrServer.scala 105:45]
  wire [66:0] _GEN_141 = {{3'd0}, rAddr}; // @[virtContAddrServer.scala 105:36]
  wire [66:0] _io_read_address_bits_T_2 = _GEN_141 + _io_read_address_bits_T; // @[virtContAddrServer.scala 105:36]
  wire [63:0] _GEN_112 = 4'h1 == burstCounter ? continuationsRegisters_1 : continuationsRegisters_0; // @[virtContAddrServer.scala 106:{27,27}]
  wire [63:0] _GEN_113 = 4'h2 == burstCounter ? continuationsRegisters_2 : _GEN_112; // @[virtContAddrServer.scala 106:{27,27}]
  wire [63:0] _GEN_114 = 4'h3 == burstCounter ? continuationsRegisters_3 : _GEN_113; // @[virtContAddrServer.scala 106:{27,27}]
  wire [63:0] _GEN_115 = 4'h4 == burstCounter ? continuationsRegisters_4 : _GEN_114; // @[virtContAddrServer.scala 106:{27,27}]
  wire [63:0] _GEN_116 = 4'h5 == burstCounter ? continuationsRegisters_5 : _GEN_115; // @[virtContAddrServer.scala 106:{27,27}]
  wire [63:0] _GEN_117 = 4'h6 == burstCounter ? continuationsRegisters_6 : _GEN_116; // @[virtContAddrServer.scala 106:{27,27}]
  wire [63:0] _GEN_118 = 4'h7 == burstCounter ? continuationsRegisters_7 : _GEN_117; // @[virtContAddrServer.scala 106:{27,27}]
  wire [63:0] _GEN_119 = 4'h8 == burstCounter ? continuationsRegisters_8 : _GEN_118; // @[virtContAddrServer.scala 106:{27,27}]
  wire [63:0] _GEN_120 = 4'h9 == burstCounter ? continuationsRegisters_9 : _GEN_119; // @[virtContAddrServer.scala 106:{27,27}]
  wire [63:0] _GEN_121 = 4'ha == burstCounter ? continuationsRegisters_10 : _GEN_120; // @[virtContAddrServer.scala 106:{27,27}]
  wire [63:0] _GEN_122 = 4'hb == burstCounter ? continuationsRegisters_11 : _GEN_121; // @[virtContAddrServer.scala 106:{27,27}]
  wire [63:0] _GEN_123 = 4'hc == burstCounter ? continuationsRegisters_12 : _GEN_122; // @[virtContAddrServer.scala 106:{27,27}]
  wire [63:0] _GEN_124 = 4'hd == burstCounter ? continuationsRegisters_13 : _GEN_123; // @[virtContAddrServer.scala 106:{27,27}]
  wire [63:0] _GEN_125 = 4'he == burstCounter ? continuationsRegisters_14 : _GEN_124; // @[virtContAddrServer.scala 106:{27,27}]
  wire [63:0] _GEN_127 = 6'h0 == rdAddr ? rPause : 64'hffffffffffffffff; // @[RegisterBlock.scala 220:10 224:38 225:16]
  wire [63:0] _GEN_128 = 6'h8 == rdAddr ? rAddr : _GEN_127; // @[RegisterBlock.scala 224:38 225:16]
  wire  _T_18 = ~reset; // @[RegisterBlock.scala 182:11]
  wire [7:0] wrReqData__bits_strb = wrReqData__deq_io_deq_bits_strb; // @[Decoupled.scala 417:19 418:14]
  wire [63:0] wrReqData__bits_data = wrReqData__deq_io_deq_bits_data; // @[Decoupled.scala 417:19 418:14]
  wire [7:0] rPause_byte_wdata = wrReqData__bits_data[7:0]; // @[Interface.scala 257:33]
  wire [7:0] rPause_byte_original = rPause[7:0]; // @[Interface.scala 258:39]
  wire [7:0] _rPause_T_8 = wrReqData__bits_strb[0] ? rPause_byte_wdata : rPause_byte_original; // @[Interface.scala 259:14]
  wire [7:0] rPause_byte_wdata_1 = wrReqData__bits_data[15:8]; // @[Interface.scala 257:33]
  wire [7:0] rPause_byte_original_1 = rPause[15:8]; // @[Interface.scala 258:39]
  wire [7:0] _rPause_T_9 = wrReqData__bits_strb[1] ? rPause_byte_wdata_1 : rPause_byte_original_1; // @[Interface.scala 259:14]
  wire [7:0] rPause_byte_wdata_2 = wrReqData__bits_data[23:16]; // @[Interface.scala 257:33]
  wire [7:0] rPause_byte_original_2 = rPause[23:16]; // @[Interface.scala 258:39]
  wire [7:0] _rPause_T_10 = wrReqData__bits_strb[2] ? rPause_byte_wdata_2 : rPause_byte_original_2; // @[Interface.scala 259:14]
  wire [7:0] rPause_byte_wdata_3 = wrReqData__bits_data[31:24]; // @[Interface.scala 257:33]
  wire [7:0] rPause_byte_original_3 = rPause[31:24]; // @[Interface.scala 258:39]
  wire [7:0] _rPause_T_11 = wrReqData__bits_strb[3] ? rPause_byte_wdata_3 : rPause_byte_original_3; // @[Interface.scala 259:14]
  wire [7:0] rPause_byte_wdata_4 = wrReqData__bits_data[39:32]; // @[Interface.scala 257:33]
  wire [7:0] rPause_byte_original_4 = rPause[39:32]; // @[Interface.scala 258:39]
  wire [7:0] _rPause_T_12 = wrReqData__bits_strb[4] ? rPause_byte_wdata_4 : rPause_byte_original_4; // @[Interface.scala 259:14]
  wire [7:0] rPause_byte_wdata_5 = wrReqData__bits_data[47:40]; // @[Interface.scala 257:33]
  wire [7:0] rPause_byte_original_5 = rPause[47:40]; // @[Interface.scala 258:39]
  wire [7:0] _rPause_T_13 = wrReqData__bits_strb[5] ? rPause_byte_wdata_5 : rPause_byte_original_5; // @[Interface.scala 259:14]
  wire [7:0] rPause_byte_wdata_6 = wrReqData__bits_data[55:48]; // @[Interface.scala 257:33]
  wire [7:0] rPause_byte_original_6 = rPause[55:48]; // @[Interface.scala 258:39]
  wire [7:0] _rPause_T_14 = wrReqData__bits_strb[6] ? rPause_byte_wdata_6 : rPause_byte_original_6; // @[Interface.scala 259:14]
  wire [7:0] rPause_byte_wdata_7 = wrReqData__bits_data[63:56]; // @[Interface.scala 257:33]
  wire [7:0] rPause_byte_original_7 = rPause[63:56]; // @[Interface.scala 258:39]
  wire [7:0] _rPause_T_15 = wrReqData__bits_strb[7] ? rPause_byte_wdata_7 : rPause_byte_original_7; // @[Interface.scala 259:14]
  wire [63:0] _rPause_T_16 = {_rPause_T_15,_rPause_T_14,_rPause_T_13,_rPause_T_12,_rPause_T_11,_rPause_T_10,_rPause_T_9,
    _rPause_T_8}; // @[Interface.scala 262:7]
  wire [7:0] rAddr_byte_original = rAddr[7:0]; // @[Interface.scala 258:39]
  wire [7:0] _rAddr_T_8 = wrReqData__bits_strb[0] ? rPause_byte_wdata : rAddr_byte_original; // @[Interface.scala 259:14]
  wire [7:0] rAddr_byte_original_1 = rAddr[15:8]; // @[Interface.scala 258:39]
  wire [7:0] _rAddr_T_9 = wrReqData__bits_strb[1] ? rPause_byte_wdata_1 : rAddr_byte_original_1; // @[Interface.scala 259:14]
  wire [7:0] rAddr_byte_original_2 = rAddr[23:16]; // @[Interface.scala 258:39]
  wire [7:0] _rAddr_T_10 = wrReqData__bits_strb[2] ? rPause_byte_wdata_2 : rAddr_byte_original_2; // @[Interface.scala 259:14]
  wire [7:0] rAddr_byte_original_3 = rAddr[31:24]; // @[Interface.scala 258:39]
  wire [7:0] _rAddr_T_11 = wrReqData__bits_strb[3] ? rPause_byte_wdata_3 : rAddr_byte_original_3; // @[Interface.scala 259:14]
  wire [7:0] rAddr_byte_original_4 = rAddr[39:32]; // @[Interface.scala 258:39]
  wire [7:0] _rAddr_T_12 = wrReqData__bits_strb[4] ? rPause_byte_wdata_4 : rAddr_byte_original_4; // @[Interface.scala 259:14]
  wire [7:0] rAddr_byte_original_5 = rAddr[47:40]; // @[Interface.scala 258:39]
  wire [7:0] _rAddr_T_13 = wrReqData__bits_strb[5] ? rPause_byte_wdata_5 : rAddr_byte_original_5; // @[Interface.scala 259:14]
  wire [7:0] rAddr_byte_original_6 = rAddr[55:48]; // @[Interface.scala 258:39]
  wire [7:0] _rAddr_T_14 = wrReqData__bits_strb[6] ? rPause_byte_wdata_6 : rAddr_byte_original_6; // @[Interface.scala 259:14]
  wire [7:0] rAddr_byte_original_7 = rAddr[63:56]; // @[Interface.scala 258:39]
  wire [7:0] _rAddr_T_15 = wrReqData__bits_strb[7] ? rPause_byte_wdata_7 : rAddr_byte_original_7; // @[Interface.scala 259:14]
  wire [63:0] _rAddr_T_16 = {_rAddr_T_15,_rAddr_T_14,_rAddr_T_13,_rAddr_T_12,_rAddr_T_11,_rAddr_T_10,_rAddr_T_9,
    _rAddr_T_8}; // @[Interface.scala 262:7]
  wire [7:0] avaialbleSize_byte_original = avaialbleSize[7:0]; // @[Interface.scala 258:39]
  wire [7:0] _avaialbleSize_T_12 = wrReqData__bits_strb[0] ? rPause_byte_wdata : avaialbleSize_byte_original; // @[Interface.scala 259:14]
  wire [7:0] avaialbleSize_byte_original_1 = avaialbleSize[15:8]; // @[Interface.scala 258:39]
  wire [7:0] _avaialbleSize_T_13 = wrReqData__bits_strb[1] ? rPause_byte_wdata_1 : avaialbleSize_byte_original_1; // @[Interface.scala 259:14]
  wire [7:0] avaialbleSize_byte_original_2 = avaialbleSize[23:16]; // @[Interface.scala 258:39]
  wire [7:0] _avaialbleSize_T_14 = wrReqData__bits_strb[2] ? rPause_byte_wdata_2 : avaialbleSize_byte_original_2; // @[Interface.scala 259:14]
  wire [7:0] avaialbleSize_byte_original_3 = avaialbleSize[31:24]; // @[Interface.scala 258:39]
  wire [7:0] _avaialbleSize_T_15 = wrReqData__bits_strb[3] ? rPause_byte_wdata_3 : avaialbleSize_byte_original_3; // @[Interface.scala 259:14]
  wire [7:0] avaialbleSize_byte_original_4 = avaialbleSize[39:32]; // @[Interface.scala 258:39]
  wire [7:0] _avaialbleSize_T_16 = wrReqData__bits_strb[4] ? rPause_byte_wdata_4 : avaialbleSize_byte_original_4; // @[Interface.scala 259:14]
  wire [7:0] avaialbleSize_byte_original_5 = avaialbleSize[47:40]; // @[Interface.scala 258:39]
  wire [7:0] _avaialbleSize_T_17 = wrReqData__bits_strb[5] ? rPause_byte_wdata_5 : avaialbleSize_byte_original_5; // @[Interface.scala 259:14]
  wire [7:0] avaialbleSize_byte_original_6 = avaialbleSize[55:48]; // @[Interface.scala 258:39]
  wire [7:0] _avaialbleSize_T_18 = wrReqData__bits_strb[6] ? rPause_byte_wdata_6 : avaialbleSize_byte_original_6; // @[Interface.scala 259:14]
  wire [7:0] avaialbleSize_byte_original_7 = avaialbleSize[63:56]; // @[Interface.scala 258:39]
  wire [7:0] _avaialbleSize_T_19 = wrReqData__bits_strb[7] ? rPause_byte_wdata_7 : avaialbleSize_byte_original_7; // @[Interface.scala 259:14]
  wire [63:0] _avaialbleSize_T_20 = {_avaialbleSize_T_19,_avaialbleSize_T_18,_avaialbleSize_T_17,_avaialbleSize_T_16,
    _avaialbleSize_T_15,_avaialbleSize_T_14,_avaialbleSize_T_13,_avaialbleSize_T_12}; // @[Interface.scala 262:7]
  Queue rdReq__deq ( // @[Decoupled.scala 377:21]
    .clock(rdReq__deq_clock),
    .reset(rdReq__deq_reset),
    .io_enq_ready(rdReq__deq_io_enq_ready),
    .io_enq_valid(rdReq__deq_io_enq_valid),
    .io_enq_bits_addr(rdReq__deq_io_enq_bits_addr),
    .io_deq_ready(rdReq__deq_io_deq_ready),
    .io_deq_valid(rdReq__deq_io_deq_valid),
    .io_deq_bits_addr(rdReq__deq_io_deq_bits_addr)
  );
  Queue wrReq__deq ( // @[Decoupled.scala 377:21]
    .clock(wrReq__deq_clock),
    .reset(wrReq__deq_reset),
    .io_enq_ready(wrReq__deq_io_enq_ready),
    .io_enq_valid(wrReq__deq_io_enq_valid),
    .io_enq_bits_addr(wrReq__deq_io_enq_bits_addr),
    .io_deq_ready(wrReq__deq_io_deq_ready),
    .io_deq_valid(wrReq__deq_io_deq_valid),
    .io_deq_bits_addr(wrReq__deq_io_deq_bits_addr)
  );
  Queue_2 wrReqData__deq ( // @[Decoupled.scala 377:21]
    .clock(wrReqData__deq_clock),
    .reset(wrReqData__deq_reset),
    .io_enq_ready(wrReqData__deq_io_enq_ready),
    .io_enq_valid(wrReqData__deq_io_enq_valid),
    .io_enq_bits_data(wrReqData__deq_io_enq_bits_data),
    .io_enq_bits_strb(wrReqData__deq_io_enq_bits_strb),
    .io_deq_ready(wrReqData__deq_io_deq_ready),
    .io_deq_valid(wrReqData__deq_io_deq_valid),
    .io_deq_bits_data(wrReqData__deq_io_deq_bits_data),
    .io_deq_bits_strb(wrReqData__deq_io_deq_bits_strb)
  );
  assign io_dataOut_valid = _T_2 ? 1'h0 : _GEN_107; // @[virtContAddrServer.scala 92:27 96:48]
  assign io_dataOut_bits = 4'hf == burstCounter ? continuationsRegisters_15 : _GEN_125; // @[virtContAddrServer.scala 106:{27,27}]
  assign io_axi_mgmt_ARREADY = rdReq__deq_io_enq_ready; // @[Decoupled.scala 381:17 RegisterBlock.scala 60:19]
  assign io_axi_mgmt_RVALID = rdReq__valid & io_axi_mgmt_RREADY; // @[RegisterBlock.scala 210:44]
  assign io_axi_mgmt_RDATA = 6'h10 == rdAddr ? avaialbleSize : _GEN_128; // @[RegisterBlock.scala 224:38 225:16]
  assign io_axi_mgmt_AWREADY = wrReq__deq_io_enq_ready; // @[Decoupled.scala 381:17 RegisterBlock.scala 60:19]
  assign io_axi_mgmt_WREADY = wrReqData__deq_io_enq_ready; // @[Decoupled.scala 381:17 RegisterBlock.scala 60:19]
  assign io_axi_mgmt_BVALID = wrReq__valid & wrReqData__valid & io_axi_mgmt_BREADY; // @[RegisterBlock.scala 241:63]
  assign io_read_address_valid = stateReg == 3'h1; // @[virtContAddrServer.scala 96:19]
  assign io_read_address_bits = _io_read_address_bits_T_2[63:0]; // @[virtContAddrServer.scala 105:27]
  assign io_read_data_ready = _T_2 ? 1'h0 : _T_3; // @[virtContAddrServer.scala 90:27 96:48]
  assign rdReq__deq_clock = clock;
  assign rdReq__deq_reset = reset;
  assign rdReq__deq_io_enq_valid = io_axi_mgmt_ARVALID; // @[RegisterBlock.scala 60:19 virtContAddrServer.scala 34:20]
  assign rdReq__deq_io_enq_bits_addr = io_axi_mgmt_ARADDR; // @[RegisterBlock.scala 60:19 virtContAddrServer.scala 34:20]
  assign rdReq__deq_io_deq_ready = rdReq__valid & io_axi_mgmt_RREADY; // @[RegisterBlock.scala 210:44]
  assign wrReq__deq_clock = clock;
  assign wrReq__deq_reset = reset;
  assign wrReq__deq_io_enq_valid = io_axi_mgmt_AWVALID; // @[RegisterBlock.scala 60:19 virtContAddrServer.scala 34:20]
  assign wrReq__deq_io_enq_bits_addr = io_axi_mgmt_AWADDR; // @[RegisterBlock.scala 60:19 virtContAddrServer.scala 34:20]
  assign wrReq__deq_io_deq_ready = wrReq__valid & wrReqData__valid & io_axi_mgmt_BREADY; // @[RegisterBlock.scala 241:63]
  assign wrReqData__deq_clock = clock;
  assign wrReqData__deq_reset = reset;
  assign wrReqData__deq_io_enq_valid = io_axi_mgmt_WVALID; // @[RegisterBlock.scala 60:19 virtContAddrServer.scala 34:20]
  assign wrReqData__deq_io_enq_bits_data = io_axi_mgmt_WDATA; // @[RegisterBlock.scala 60:19 virtContAddrServer.scala 34:20]
  assign wrReqData__deq_io_enq_bits_strb = io_axi_mgmt_WSTRB; // @[RegisterBlock.scala 60:19 virtContAddrServer.scala 34:20]
  assign wrReqData__deq_io_deq_ready = wrReq__valid & wrReqData__valid & io_axi_mgmt_BREADY; // @[RegisterBlock.scala 241:63]
  always @(posedge clock) begin
    if (reset) begin // @[virtContAddrServer.scala 37:49]
      rAddr <= 64'h0; // @[virtContAddrServer.scala 37:49]
    end else if (wrReq) begin // @[virtContAddrServer.scala 113:27]
      if (6'h8 == wrAddr) begin // @[RegisterBlock.scala 252:38]
        rAddr <= _rAddr_T_16; // @[RegisterBlock.scala 118:11]
      end
    end
    if (reset) begin // @[virtContAddrServer.scala 38:49]
      rPause <= 64'h0; // @[virtContAddrServer.scala 38:49]
    end else if (wrReq) begin // @[virtContAddrServer.scala 113:27]
      if (6'h0 == wrAddr) begin // @[RegisterBlock.scala 252:38]
        rPause <= _rPause_T_16; // @[RegisterBlock.scala 118:11]
      end else begin
        rPause <= _GEN_86;
      end
    end else begin
      rPause <= _GEN_86;
    end
    if (reset) begin // @[virtContAddrServer.scala 39:49]
      avaialbleSize <= 64'h0; // @[virtContAddrServer.scala 39:49]
    end else if (wrReq) begin // @[virtContAddrServer.scala 113:27]
      if (6'h10 == wrAddr) begin // @[RegisterBlock.scala 252:38]
        avaialbleSize <= _avaialbleSize_T_20; // @[RegisterBlock.scala 118:11]
      end else begin
        avaialbleSize <= _GEN_104;
      end
    end else begin
      avaialbleSize <= _GEN_104;
    end
    if (reset) begin // @[virtContAddrServer.scala 40:49]
      stateReg <= 3'h0; // @[virtContAddrServer.scala 40:49]
    end else if (stateReg == 3'h0) begin // @[virtContAddrServer.scala 51:34]
      if (avaialbleSize >= 64'h10) begin // @[virtContAddrServer.scala 52:52]
        stateReg <= 3'h1; // @[virtContAddrServer.scala 53:22]
      end else begin
        stateReg <= 3'h4; // @[virtContAddrServer.scala 55:22]
      end
    end else if (stateReg == 3'h1) begin // @[virtContAddrServer.scala 58:54]
      if (io_read_address_ready) begin // @[virtContAddrServer.scala 59:36]
        stateReg <= 3'h2; // @[virtContAddrServer.scala 60:26]
      end
    end else if (stateReg == 3'h2) begin // @[virtContAddrServer.scala 63:44]
      stateReg <= _GEN_38;
    end else begin
      stateReg <= _GEN_46;
    end
    if (reset) begin // @[virtContAddrServer.scala 43:49]
      continuationsRegisters_0 <= 64'h0; // @[virtContAddrServer.scala 43:49]
    end else if (!(stateReg == 3'h0)) begin // @[virtContAddrServer.scala 51:34]
      if (!(stateReg == 3'h1)) begin // @[virtContAddrServer.scala 58:54]
        if (stateReg == 3'h2) begin // @[virtContAddrServer.scala 63:44]
          continuationsRegisters_0 <= _GEN_20;
        end
      end
    end
    if (reset) begin // @[virtContAddrServer.scala 43:49]
      continuationsRegisters_1 <= 64'h0; // @[virtContAddrServer.scala 43:49]
    end else if (!(stateReg == 3'h0)) begin // @[virtContAddrServer.scala 51:34]
      if (!(stateReg == 3'h1)) begin // @[virtContAddrServer.scala 58:54]
        if (stateReg == 3'h2) begin // @[virtContAddrServer.scala 63:44]
          continuationsRegisters_1 <= _GEN_21;
        end
      end
    end
    if (reset) begin // @[virtContAddrServer.scala 43:49]
      continuationsRegisters_2 <= 64'h0; // @[virtContAddrServer.scala 43:49]
    end else if (!(stateReg == 3'h0)) begin // @[virtContAddrServer.scala 51:34]
      if (!(stateReg == 3'h1)) begin // @[virtContAddrServer.scala 58:54]
        if (stateReg == 3'h2) begin // @[virtContAddrServer.scala 63:44]
          continuationsRegisters_2 <= _GEN_22;
        end
      end
    end
    if (reset) begin // @[virtContAddrServer.scala 43:49]
      continuationsRegisters_3 <= 64'h0; // @[virtContAddrServer.scala 43:49]
    end else if (!(stateReg == 3'h0)) begin // @[virtContAddrServer.scala 51:34]
      if (!(stateReg == 3'h1)) begin // @[virtContAddrServer.scala 58:54]
        if (stateReg == 3'h2) begin // @[virtContAddrServer.scala 63:44]
          continuationsRegisters_3 <= _GEN_23;
        end
      end
    end
    if (reset) begin // @[virtContAddrServer.scala 43:49]
      continuationsRegisters_4 <= 64'h0; // @[virtContAddrServer.scala 43:49]
    end else if (!(stateReg == 3'h0)) begin // @[virtContAddrServer.scala 51:34]
      if (!(stateReg == 3'h1)) begin // @[virtContAddrServer.scala 58:54]
        if (stateReg == 3'h2) begin // @[virtContAddrServer.scala 63:44]
          continuationsRegisters_4 <= _GEN_24;
        end
      end
    end
    if (reset) begin // @[virtContAddrServer.scala 43:49]
      continuationsRegisters_5 <= 64'h0; // @[virtContAddrServer.scala 43:49]
    end else if (!(stateReg == 3'h0)) begin // @[virtContAddrServer.scala 51:34]
      if (!(stateReg == 3'h1)) begin // @[virtContAddrServer.scala 58:54]
        if (stateReg == 3'h2) begin // @[virtContAddrServer.scala 63:44]
          continuationsRegisters_5 <= _GEN_25;
        end
      end
    end
    if (reset) begin // @[virtContAddrServer.scala 43:49]
      continuationsRegisters_6 <= 64'h0; // @[virtContAddrServer.scala 43:49]
    end else if (!(stateReg == 3'h0)) begin // @[virtContAddrServer.scala 51:34]
      if (!(stateReg == 3'h1)) begin // @[virtContAddrServer.scala 58:54]
        if (stateReg == 3'h2) begin // @[virtContAddrServer.scala 63:44]
          continuationsRegisters_6 <= _GEN_26;
        end
      end
    end
    if (reset) begin // @[virtContAddrServer.scala 43:49]
      continuationsRegisters_7 <= 64'h0; // @[virtContAddrServer.scala 43:49]
    end else if (!(stateReg == 3'h0)) begin // @[virtContAddrServer.scala 51:34]
      if (!(stateReg == 3'h1)) begin // @[virtContAddrServer.scala 58:54]
        if (stateReg == 3'h2) begin // @[virtContAddrServer.scala 63:44]
          continuationsRegisters_7 <= _GEN_27;
        end
      end
    end
    if (reset) begin // @[virtContAddrServer.scala 43:49]
      continuationsRegisters_8 <= 64'h0; // @[virtContAddrServer.scala 43:49]
    end else if (!(stateReg == 3'h0)) begin // @[virtContAddrServer.scala 51:34]
      if (!(stateReg == 3'h1)) begin // @[virtContAddrServer.scala 58:54]
        if (stateReg == 3'h2) begin // @[virtContAddrServer.scala 63:44]
          continuationsRegisters_8 <= _GEN_28;
        end
      end
    end
    if (reset) begin // @[virtContAddrServer.scala 43:49]
      continuationsRegisters_9 <= 64'h0; // @[virtContAddrServer.scala 43:49]
    end else if (!(stateReg == 3'h0)) begin // @[virtContAddrServer.scala 51:34]
      if (!(stateReg == 3'h1)) begin // @[virtContAddrServer.scala 58:54]
        if (stateReg == 3'h2) begin // @[virtContAddrServer.scala 63:44]
          continuationsRegisters_9 <= _GEN_29;
        end
      end
    end
    if (reset) begin // @[virtContAddrServer.scala 43:49]
      continuationsRegisters_10 <= 64'h0; // @[virtContAddrServer.scala 43:49]
    end else if (!(stateReg == 3'h0)) begin // @[virtContAddrServer.scala 51:34]
      if (!(stateReg == 3'h1)) begin // @[virtContAddrServer.scala 58:54]
        if (stateReg == 3'h2) begin // @[virtContAddrServer.scala 63:44]
          continuationsRegisters_10 <= _GEN_30;
        end
      end
    end
    if (reset) begin // @[virtContAddrServer.scala 43:49]
      continuationsRegisters_11 <= 64'h0; // @[virtContAddrServer.scala 43:49]
    end else if (!(stateReg == 3'h0)) begin // @[virtContAddrServer.scala 51:34]
      if (!(stateReg == 3'h1)) begin // @[virtContAddrServer.scala 58:54]
        if (stateReg == 3'h2) begin // @[virtContAddrServer.scala 63:44]
          continuationsRegisters_11 <= _GEN_31;
        end
      end
    end
    if (reset) begin // @[virtContAddrServer.scala 43:49]
      continuationsRegisters_12 <= 64'h0; // @[virtContAddrServer.scala 43:49]
    end else if (!(stateReg == 3'h0)) begin // @[virtContAddrServer.scala 51:34]
      if (!(stateReg == 3'h1)) begin // @[virtContAddrServer.scala 58:54]
        if (stateReg == 3'h2) begin // @[virtContAddrServer.scala 63:44]
          continuationsRegisters_12 <= _GEN_32;
        end
      end
    end
    if (reset) begin // @[virtContAddrServer.scala 43:49]
      continuationsRegisters_13 <= 64'h0; // @[virtContAddrServer.scala 43:49]
    end else if (!(stateReg == 3'h0)) begin // @[virtContAddrServer.scala 51:34]
      if (!(stateReg == 3'h1)) begin // @[virtContAddrServer.scala 58:54]
        if (stateReg == 3'h2) begin // @[virtContAddrServer.scala 63:44]
          continuationsRegisters_13 <= _GEN_33;
        end
      end
    end
    if (reset) begin // @[virtContAddrServer.scala 43:49]
      continuationsRegisters_14 <= 64'h0; // @[virtContAddrServer.scala 43:49]
    end else if (!(stateReg == 3'h0)) begin // @[virtContAddrServer.scala 51:34]
      if (!(stateReg == 3'h1)) begin // @[virtContAddrServer.scala 58:54]
        if (stateReg == 3'h2) begin // @[virtContAddrServer.scala 63:44]
          continuationsRegisters_14 <= _GEN_34;
        end
      end
    end
    if (reset) begin // @[virtContAddrServer.scala 43:49]
      continuationsRegisters_15 <= 64'h0; // @[virtContAddrServer.scala 43:49]
    end else if (!(stateReg == 3'h0)) begin // @[virtContAddrServer.scala 51:34]
      if (!(stateReg == 3'h1)) begin // @[virtContAddrServer.scala 58:54]
        if (stateReg == 3'h2) begin // @[virtContAddrServer.scala 63:44]
          continuationsRegisters_15 <= _GEN_35;
        end
      end
    end
    if (reset) begin // @[virtContAddrServer.scala 44:49]
      burstCounter <= 4'hf; // @[virtContAddrServer.scala 44:49]
    end else if (!(stateReg == 3'h0)) begin // @[virtContAddrServer.scala 51:34]
      if (stateReg == 3'h1) begin // @[virtContAddrServer.scala 58:54]
        if (io_read_address_ready) begin // @[virtContAddrServer.scala 59:36]
          burstCounter <= 4'hf; // @[virtContAddrServer.scala 61:26]
        end
      end else if (stateReg == 3'h2) begin // @[virtContAddrServer.scala 63:44]
        burstCounter <= _GEN_40;
      end else begin
        burstCounter <= _GEN_45;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (rdReq & ~reset & ~rdReq) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegisterBlock.scala:182 assert(rdReq)\n"); // @[RegisterBlock.scala 182:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~rdReq & (rdReq & ~reset)) begin
          $fatal; // @[RegisterBlock.scala 182:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (wrReq & _T_18 & ~wrReq) begin
          $fwrite(32'h80000002,"Assertion failed\n    at RegisterBlock.scala:198 assert(wrReq)\n"); // @[RegisterBlock.scala 198:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~wrReq & (wrReq & _T_18)) begin
          $fatal; // @[RegisterBlock.scala 198:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  rAddr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  rPause = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  avaialbleSize = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  stateReg = _RAND_3[2:0];
  _RAND_4 = {2{`RANDOM}};
  continuationsRegisters_0 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  continuationsRegisters_1 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  continuationsRegisters_2 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  continuationsRegisters_3 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  continuationsRegisters_4 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  continuationsRegisters_5 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  continuationsRegisters_6 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  continuationsRegisters_7 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  continuationsRegisters_8 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  continuationsRegisters_9 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  continuationsRegisters_10 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  continuationsRegisters_11 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  continuationsRegisters_12 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  continuationsRegisters_13 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  continuationsRegisters_14 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  continuationsRegisters_15 = _RAND_19[63:0];
  _RAND_20 = {1{`RANDOM}};
  burstCounter = _RAND_20[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module readyValidMem_1(
  output        io_read_address_ready,
  input         io_read_address_valid,
  input  [63:0] io_read_address_bits,
  input         io_read_data_ready,
  output        io_read_data_valid,
  output [63:0] io_read_data_bits,
  input         axi_ARREADY,
  output        axi_ARVALID,
  output [63:0] axi_ARADDR,
  output        axi_RREADY,
  input         axi_RVALID,
  input  [63:0] axi_RDATA
);
  assign io_read_address_ready = axi_ARREADY; // @[readyValidMem.scala 155:31]
  assign io_read_data_valid = axi_RVALID; // @[readyValidMem.scala 171:31]
  assign io_read_data_bits = axi_RDATA; // @[readyValidMem.scala 172:31]
  assign axi_ARVALID = io_read_address_valid; // @[readyValidMem.scala 153:31]
  assign axi_ARADDR = io_read_address_bits; // @[readyValidMem.scala 154:31]
  assign axi_RREADY = io_read_data_ready; // @[readyValidMem.scala 169:31]
endmodule
module continuationAllocationSide(
  input         clock,
  input         reset,
  input         io_contOut_0_TREADY,
  output        io_contOut_0_TVALID,
  output [63:0] io_contOut_0_TDATA,
  input         io_contOut_1_TREADY,
  output        io_contOut_1_TVALID,
  output [63:0] io_contOut_1_TDATA,
  input         io_contOut_2_TREADY,
  output        io_contOut_2_TVALID,
  output [63:0] io_contOut_2_TDATA,
  input         io_contOut_3_TREADY,
  output        io_contOut_3_TVALID,
  output [63:0] io_contOut_3_TDATA,
  input         io_contOut_4_TREADY,
  output        io_contOut_4_TVALID,
  output [63:0] io_contOut_4_TDATA,
  input         io_contOut_5_TREADY,
  output        io_contOut_5_TVALID,
  output [63:0] io_contOut_5_TDATA,
  input         io_contOut_6_TREADY,
  output        io_contOut_6_TVALID,
  output [63:0] io_contOut_6_TDATA,
  input         io_contOut_7_TREADY,
  output        io_contOut_7_TVALID,
  output [63:0] io_contOut_7_TDATA,
  input         io_contOut_8_TREADY,
  output        io_contOut_8_TVALID,
  output [63:0] io_contOut_8_TDATA,
  input         io_contOut_9_TREADY,
  output        io_contOut_9_TVALID,
  output [63:0] io_contOut_9_TDATA,
  input         io_contOut_10_TREADY,
  output        io_contOut_10_TVALID,
  output [63:0] io_contOut_10_TDATA,
  input         io_contOut_11_TREADY,
  output        io_contOut_11_TVALID,
  output [63:0] io_contOut_11_TDATA,
  input         io_contOut_12_TREADY,
  output        io_contOut_12_TVALID,
  output [63:0] io_contOut_12_TDATA,
  input         io_contOut_13_TREADY,
  output        io_contOut_13_TVALID,
  output [63:0] io_contOut_13_TDATA,
  input         io_contOut_14_TREADY,
  output        io_contOut_14_TVALID,
  output [63:0] io_contOut_14_TDATA,
  input         io_contOut_15_TREADY,
  output        io_contOut_15_TVALID,
  output [63:0] io_contOut_15_TDATA,
  input         io_contOut_16_TREADY,
  output        io_contOut_16_TVALID,
  output [63:0] io_contOut_16_TDATA,
  input         io_contOut_17_TREADY,
  output        io_contOut_17_TVALID,
  output [63:0] io_contOut_17_TDATA,
  input         io_contOut_18_TREADY,
  output        io_contOut_18_TVALID,
  output [63:0] io_contOut_18_TDATA,
  input         io_contOut_19_TREADY,
  output        io_contOut_19_TVALID,
  output [63:0] io_contOut_19_TDATA,
  input         io_contOut_20_TREADY,
  output        io_contOut_20_TVALID,
  output [63:0] io_contOut_20_TDATA,
  input         io_contOut_21_TREADY,
  output        io_contOut_21_TVALID,
  output [63:0] io_contOut_21_TDATA,
  input         io_contOut_22_TREADY,
  output        io_contOut_22_TVALID,
  output [63:0] io_contOut_22_TDATA,
  input         io_contOut_23_TREADY,
  output        io_contOut_23_TVALID,
  output [63:0] io_contOut_23_TDATA,
  input         io_contOut_24_TREADY,
  output        io_contOut_24_TVALID,
  output [63:0] io_contOut_24_TDATA,
  input         io_contOut_25_TREADY,
  output        io_contOut_25_TVALID,
  output [63:0] io_contOut_25_TDATA,
  input         io_contOut_26_TREADY,
  output        io_contOut_26_TVALID,
  output [63:0] io_contOut_26_TDATA,
  input         io_contOut_27_TREADY,
  output        io_contOut_27_TVALID,
  output [63:0] io_contOut_27_TDATA,
  input         io_contOut_28_TREADY,
  output        io_contOut_28_TVALID,
  output [63:0] io_contOut_28_TDATA,
  input         io_contOut_29_TREADY,
  output        io_contOut_29_TVALID,
  output [63:0] io_contOut_29_TDATA,
  input         io_contOut_30_TREADY,
  output        io_contOut_30_TVALID,
  output [63:0] io_contOut_30_TDATA,
  input         io_contOut_31_TREADY,
  output        io_contOut_31_TVALID,
  output [63:0] io_contOut_31_TDATA,
  input         io_contOut_32_TREADY,
  output        io_contOut_32_TVALID,
  output [63:0] io_contOut_32_TDATA,
  input         io_contOut_33_TREADY,
  output        io_contOut_33_TVALID,
  output [63:0] io_contOut_33_TDATA,
  input         io_contOut_34_TREADY,
  output        io_contOut_34_TVALID,
  output [63:0] io_contOut_34_TDATA,
  input         io_contOut_35_TREADY,
  output        io_contOut_35_TVALID,
  output [63:0] io_contOut_35_TDATA,
  input         io_contOut_36_TREADY,
  output        io_contOut_36_TVALID,
  output [63:0] io_contOut_36_TDATA,
  input         io_contOut_37_TREADY,
  output        io_contOut_37_TVALID,
  output [63:0] io_contOut_37_TDATA,
  input         io_contOut_38_TREADY,
  output        io_contOut_38_TVALID,
  output [63:0] io_contOut_38_TDATA,
  input         io_contOut_39_TREADY,
  output        io_contOut_39_TVALID,
  output [63:0] io_contOut_39_TDATA,
  input         io_contOut_40_TREADY,
  output        io_contOut_40_TVALID,
  output [63:0] io_contOut_40_TDATA,
  input         io_contOut_41_TREADY,
  output        io_contOut_41_TVALID,
  output [63:0] io_contOut_41_TDATA,
  input         io_contOut_42_TREADY,
  output        io_contOut_42_TVALID,
  output [63:0] io_contOut_42_TDATA,
  input         io_contOut_43_TREADY,
  output        io_contOut_43_TVALID,
  output [63:0] io_contOut_43_TDATA,
  input         io_contOut_44_TREADY,
  output        io_contOut_44_TVALID,
  output [63:0] io_contOut_44_TDATA,
  input         io_contOut_45_TREADY,
  output        io_contOut_45_TVALID,
  output [63:0] io_contOut_45_TDATA,
  input         io_contOut_46_TREADY,
  output        io_contOut_46_TVALID,
  output [63:0] io_contOut_46_TDATA,
  input         io_contOut_47_TREADY,
  output        io_contOut_47_TVALID,
  output [63:0] io_contOut_47_TDATA,
  input         io_contOut_48_TREADY,
  output        io_contOut_48_TVALID,
  output [63:0] io_contOut_48_TDATA,
  input         io_contOut_49_TREADY,
  output        io_contOut_49_TVALID,
  output [63:0] io_contOut_49_TDATA,
  input         io_contOut_50_TREADY,
  output        io_contOut_50_TVALID,
  output [63:0] io_contOut_50_TDATA,
  input         io_contOut_51_TREADY,
  output        io_contOut_51_TVALID,
  output [63:0] io_contOut_51_TDATA,
  input         io_contOut_52_TREADY,
  output        io_contOut_52_TVALID,
  output [63:0] io_contOut_52_TDATA,
  input         io_contOut_53_TREADY,
  output        io_contOut_53_TVALID,
  output [63:0] io_contOut_53_TDATA,
  input         io_contOut_54_TREADY,
  output        io_contOut_54_TVALID,
  output [63:0] io_contOut_54_TDATA,
  input         io_contOut_55_TREADY,
  output        io_contOut_55_TVALID,
  output [63:0] io_contOut_55_TDATA,
  input         io_contOut_56_TREADY,
  output        io_contOut_56_TVALID,
  output [63:0] io_contOut_56_TDATA,
  input         io_contOut_57_TREADY,
  output        io_contOut_57_TVALID,
  output [63:0] io_contOut_57_TDATA,
  input         io_contOut_58_TREADY,
  output        io_contOut_58_TVALID,
  output [63:0] io_contOut_58_TDATA,
  input         io_contOut_59_TREADY,
  output        io_contOut_59_TVALID,
  output [63:0] io_contOut_59_TDATA,
  input         io_contOut_60_TREADY,
  output        io_contOut_60_TVALID,
  output [63:0] io_contOut_60_TDATA,
  input         io_contOut_61_TREADY,
  output        io_contOut_61_TVALID,
  output [63:0] io_contOut_61_TDATA,
  input         io_contOut_62_TREADY,
  output        io_contOut_62_TVALID,
  output [63:0] io_contOut_62_TDATA,
  input         io_contOut_63_TREADY,
  output        io_contOut_63_TVALID,
  output [63:0] io_contOut_63_TDATA,
  output        io_axi_mgmt_vcas_0_ARREADY,
  input         io_axi_mgmt_vcas_0_ARVALID,
  input  [5:0]  io_axi_mgmt_vcas_0_ARADDR,
  input         io_axi_mgmt_vcas_0_RREADY,
  output        io_axi_mgmt_vcas_0_RVALID,
  output [63:0] io_axi_mgmt_vcas_0_RDATA,
  output        io_axi_mgmt_vcas_0_AWREADY,
  input         io_axi_mgmt_vcas_0_AWVALID,
  input  [5:0]  io_axi_mgmt_vcas_0_AWADDR,
  output        io_axi_mgmt_vcas_0_WREADY,
  input         io_axi_mgmt_vcas_0_WVALID,
  input  [63:0] io_axi_mgmt_vcas_0_WDATA,
  input  [7:0]  io_axi_mgmt_vcas_0_WSTRB,
  input         io_axi_mgmt_vcas_0_BREADY,
  output        io_axi_mgmt_vcas_0_BVALID,
  input         io_vcas_axi_full_0_ARREADY,
  output        io_vcas_axi_full_0_ARVALID,
  output [63:0] io_vcas_axi_full_0_ARADDR,
  output        io_vcas_axi_full_0_RREADY,
  input         io_vcas_axi_full_0_RVALID,
  input  [63:0] io_vcas_axi_full_0_RDATA
);
  wire  continuationNetwork_clock; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_reset; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connVCAS_0_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connVCAS_0_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connVCAS_0_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_0_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_0_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_0_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_1_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_1_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_1_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_2_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_2_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_2_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_3_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_3_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_3_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_4_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_4_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_4_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_5_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_5_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_5_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_6_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_6_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_6_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_7_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_7_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_7_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_8_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_8_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_8_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_9_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_9_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_9_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_10_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_10_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_10_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_11_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_11_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_11_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_12_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_12_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_12_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_13_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_13_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_13_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_14_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_14_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_14_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_15_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_15_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_15_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_16_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_16_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_16_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_17_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_17_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_17_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_18_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_18_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_18_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_19_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_19_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_19_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_20_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_20_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_20_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_21_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_21_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_21_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_22_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_22_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_22_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_23_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_23_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_23_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_24_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_24_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_24_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_25_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_25_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_25_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_26_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_26_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_26_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_27_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_27_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_27_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_28_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_28_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_28_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_29_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_29_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_29_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_30_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_30_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_30_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_31_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_31_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_31_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_32_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_32_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_32_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_33_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_33_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_33_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_34_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_34_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_34_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_35_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_35_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_35_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_36_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_36_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_36_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_37_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_37_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_37_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_38_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_38_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_38_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_39_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_39_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_39_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_40_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_40_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_40_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_41_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_41_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_41_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_42_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_42_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_42_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_43_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_43_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_43_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_44_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_44_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_44_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_45_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_45_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_45_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_46_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_46_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_46_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_47_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_47_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_47_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_48_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_48_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_48_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_49_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_49_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_49_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_50_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_50_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_50_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_51_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_51_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_51_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_52_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_52_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_52_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_53_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_53_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_53_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_54_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_54_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_54_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_55_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_55_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_55_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_56_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_56_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_56_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_57_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_57_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_57_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_58_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_58_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_58_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_59_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_59_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_59_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_60_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_60_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_60_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_61_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_61_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_61_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_62_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_62_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_62_bits; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_63_ready; // @[continuationAllocationSide.scala 52:37]
  wire  continuationNetwork_io_connPE_63_valid; // @[continuationAllocationSide.scala 52:37]
  wire [63:0] continuationNetwork_io_connPE_63_bits; // @[continuationAllocationSide.scala 52:37]
  wire  vcas_0_clock; // @[continuationAllocationSide.scala 58:42]
  wire  vcas_0_reset; // @[continuationAllocationSide.scala 58:42]
  wire  vcas_0_io_dataOut_ready; // @[continuationAllocationSide.scala 58:42]
  wire  vcas_0_io_dataOut_valid; // @[continuationAllocationSide.scala 58:42]
  wire [63:0] vcas_0_io_dataOut_bits; // @[continuationAllocationSide.scala 58:42]
  wire  vcas_0_io_axi_mgmt_ARREADY; // @[continuationAllocationSide.scala 58:42]
  wire  vcas_0_io_axi_mgmt_ARVALID; // @[continuationAllocationSide.scala 58:42]
  wire [5:0] vcas_0_io_axi_mgmt_ARADDR; // @[continuationAllocationSide.scala 58:42]
  wire  vcas_0_io_axi_mgmt_RREADY; // @[continuationAllocationSide.scala 58:42]
  wire  vcas_0_io_axi_mgmt_RVALID; // @[continuationAllocationSide.scala 58:42]
  wire [63:0] vcas_0_io_axi_mgmt_RDATA; // @[continuationAllocationSide.scala 58:42]
  wire  vcas_0_io_axi_mgmt_AWREADY; // @[continuationAllocationSide.scala 58:42]
  wire  vcas_0_io_axi_mgmt_AWVALID; // @[continuationAllocationSide.scala 58:42]
  wire [5:0] vcas_0_io_axi_mgmt_AWADDR; // @[continuationAllocationSide.scala 58:42]
  wire  vcas_0_io_axi_mgmt_WREADY; // @[continuationAllocationSide.scala 58:42]
  wire  vcas_0_io_axi_mgmt_WVALID; // @[continuationAllocationSide.scala 58:42]
  wire [63:0] vcas_0_io_axi_mgmt_WDATA; // @[continuationAllocationSide.scala 58:42]
  wire [7:0] vcas_0_io_axi_mgmt_WSTRB; // @[continuationAllocationSide.scala 58:42]
  wire  vcas_0_io_axi_mgmt_BREADY; // @[continuationAllocationSide.scala 58:42]
  wire  vcas_0_io_axi_mgmt_BVALID; // @[continuationAllocationSide.scala 58:42]
  wire  vcas_0_io_read_address_ready; // @[continuationAllocationSide.scala 58:42]
  wire  vcas_0_io_read_address_valid; // @[continuationAllocationSide.scala 58:42]
  wire [63:0] vcas_0_io_read_address_bits; // @[continuationAllocationSide.scala 58:42]
  wire  vcas_0_io_read_data_ready; // @[continuationAllocationSide.scala 58:42]
  wire  vcas_0_io_read_data_valid; // @[continuationAllocationSide.scala 58:42]
  wire [63:0] vcas_0_io_read_data_bits; // @[continuationAllocationSide.scala 58:42]
  wire  vcasRvmRO_0_io_read_address_ready; // @[continuationAllocationSide.scala 71:47]
  wire  vcasRvmRO_0_io_read_address_valid; // @[continuationAllocationSide.scala 71:47]
  wire [63:0] vcasRvmRO_0_io_read_address_bits; // @[continuationAllocationSide.scala 71:47]
  wire  vcasRvmRO_0_io_read_data_ready; // @[continuationAllocationSide.scala 71:47]
  wire  vcasRvmRO_0_io_read_data_valid; // @[continuationAllocationSide.scala 71:47]
  wire [63:0] vcasRvmRO_0_io_read_data_bits; // @[continuationAllocationSide.scala 71:47]
  wire  vcasRvmRO_0_axi_ARREADY; // @[continuationAllocationSide.scala 71:47]
  wire  vcasRvmRO_0_axi_ARVALID; // @[continuationAllocationSide.scala 71:47]
  wire [63:0] vcasRvmRO_0_axi_ARADDR; // @[continuationAllocationSide.scala 71:47]
  wire  vcasRvmRO_0_axi_RREADY; // @[continuationAllocationSide.scala 71:47]
  wire  vcasRvmRO_0_axi_RVALID; // @[continuationAllocationSide.scala 71:47]
  wire [63:0] vcasRvmRO_0_axi_RDATA; // @[continuationAllocationSide.scala 71:47]
  contNetwork continuationNetwork ( // @[continuationAllocationSide.scala 52:37]
    .clock(continuationNetwork_clock),
    .reset(continuationNetwork_reset),
    .io_connVCAS_0_ready(continuationNetwork_io_connVCAS_0_ready),
    .io_connVCAS_0_valid(continuationNetwork_io_connVCAS_0_valid),
    .io_connVCAS_0_bits(continuationNetwork_io_connVCAS_0_bits),
    .io_connPE_0_ready(continuationNetwork_io_connPE_0_ready),
    .io_connPE_0_valid(continuationNetwork_io_connPE_0_valid),
    .io_connPE_0_bits(continuationNetwork_io_connPE_0_bits),
    .io_connPE_1_ready(continuationNetwork_io_connPE_1_ready),
    .io_connPE_1_valid(continuationNetwork_io_connPE_1_valid),
    .io_connPE_1_bits(continuationNetwork_io_connPE_1_bits),
    .io_connPE_2_ready(continuationNetwork_io_connPE_2_ready),
    .io_connPE_2_valid(continuationNetwork_io_connPE_2_valid),
    .io_connPE_2_bits(continuationNetwork_io_connPE_2_bits),
    .io_connPE_3_ready(continuationNetwork_io_connPE_3_ready),
    .io_connPE_3_valid(continuationNetwork_io_connPE_3_valid),
    .io_connPE_3_bits(continuationNetwork_io_connPE_3_bits),
    .io_connPE_4_ready(continuationNetwork_io_connPE_4_ready),
    .io_connPE_4_valid(continuationNetwork_io_connPE_4_valid),
    .io_connPE_4_bits(continuationNetwork_io_connPE_4_bits),
    .io_connPE_5_ready(continuationNetwork_io_connPE_5_ready),
    .io_connPE_5_valid(continuationNetwork_io_connPE_5_valid),
    .io_connPE_5_bits(continuationNetwork_io_connPE_5_bits),
    .io_connPE_6_ready(continuationNetwork_io_connPE_6_ready),
    .io_connPE_6_valid(continuationNetwork_io_connPE_6_valid),
    .io_connPE_6_bits(continuationNetwork_io_connPE_6_bits),
    .io_connPE_7_ready(continuationNetwork_io_connPE_7_ready),
    .io_connPE_7_valid(continuationNetwork_io_connPE_7_valid),
    .io_connPE_7_bits(continuationNetwork_io_connPE_7_bits),
    .io_connPE_8_ready(continuationNetwork_io_connPE_8_ready),
    .io_connPE_8_valid(continuationNetwork_io_connPE_8_valid),
    .io_connPE_8_bits(continuationNetwork_io_connPE_8_bits),
    .io_connPE_9_ready(continuationNetwork_io_connPE_9_ready),
    .io_connPE_9_valid(continuationNetwork_io_connPE_9_valid),
    .io_connPE_9_bits(continuationNetwork_io_connPE_9_bits),
    .io_connPE_10_ready(continuationNetwork_io_connPE_10_ready),
    .io_connPE_10_valid(continuationNetwork_io_connPE_10_valid),
    .io_connPE_10_bits(continuationNetwork_io_connPE_10_bits),
    .io_connPE_11_ready(continuationNetwork_io_connPE_11_ready),
    .io_connPE_11_valid(continuationNetwork_io_connPE_11_valid),
    .io_connPE_11_bits(continuationNetwork_io_connPE_11_bits),
    .io_connPE_12_ready(continuationNetwork_io_connPE_12_ready),
    .io_connPE_12_valid(continuationNetwork_io_connPE_12_valid),
    .io_connPE_12_bits(continuationNetwork_io_connPE_12_bits),
    .io_connPE_13_ready(continuationNetwork_io_connPE_13_ready),
    .io_connPE_13_valid(continuationNetwork_io_connPE_13_valid),
    .io_connPE_13_bits(continuationNetwork_io_connPE_13_bits),
    .io_connPE_14_ready(continuationNetwork_io_connPE_14_ready),
    .io_connPE_14_valid(continuationNetwork_io_connPE_14_valid),
    .io_connPE_14_bits(continuationNetwork_io_connPE_14_bits),
    .io_connPE_15_ready(continuationNetwork_io_connPE_15_ready),
    .io_connPE_15_valid(continuationNetwork_io_connPE_15_valid),
    .io_connPE_15_bits(continuationNetwork_io_connPE_15_bits),
    .io_connPE_16_ready(continuationNetwork_io_connPE_16_ready),
    .io_connPE_16_valid(continuationNetwork_io_connPE_16_valid),
    .io_connPE_16_bits(continuationNetwork_io_connPE_16_bits),
    .io_connPE_17_ready(continuationNetwork_io_connPE_17_ready),
    .io_connPE_17_valid(continuationNetwork_io_connPE_17_valid),
    .io_connPE_17_bits(continuationNetwork_io_connPE_17_bits),
    .io_connPE_18_ready(continuationNetwork_io_connPE_18_ready),
    .io_connPE_18_valid(continuationNetwork_io_connPE_18_valid),
    .io_connPE_18_bits(continuationNetwork_io_connPE_18_bits),
    .io_connPE_19_ready(continuationNetwork_io_connPE_19_ready),
    .io_connPE_19_valid(continuationNetwork_io_connPE_19_valid),
    .io_connPE_19_bits(continuationNetwork_io_connPE_19_bits),
    .io_connPE_20_ready(continuationNetwork_io_connPE_20_ready),
    .io_connPE_20_valid(continuationNetwork_io_connPE_20_valid),
    .io_connPE_20_bits(continuationNetwork_io_connPE_20_bits),
    .io_connPE_21_ready(continuationNetwork_io_connPE_21_ready),
    .io_connPE_21_valid(continuationNetwork_io_connPE_21_valid),
    .io_connPE_21_bits(continuationNetwork_io_connPE_21_bits),
    .io_connPE_22_ready(continuationNetwork_io_connPE_22_ready),
    .io_connPE_22_valid(continuationNetwork_io_connPE_22_valid),
    .io_connPE_22_bits(continuationNetwork_io_connPE_22_bits),
    .io_connPE_23_ready(continuationNetwork_io_connPE_23_ready),
    .io_connPE_23_valid(continuationNetwork_io_connPE_23_valid),
    .io_connPE_23_bits(continuationNetwork_io_connPE_23_bits),
    .io_connPE_24_ready(continuationNetwork_io_connPE_24_ready),
    .io_connPE_24_valid(continuationNetwork_io_connPE_24_valid),
    .io_connPE_24_bits(continuationNetwork_io_connPE_24_bits),
    .io_connPE_25_ready(continuationNetwork_io_connPE_25_ready),
    .io_connPE_25_valid(continuationNetwork_io_connPE_25_valid),
    .io_connPE_25_bits(continuationNetwork_io_connPE_25_bits),
    .io_connPE_26_ready(continuationNetwork_io_connPE_26_ready),
    .io_connPE_26_valid(continuationNetwork_io_connPE_26_valid),
    .io_connPE_26_bits(continuationNetwork_io_connPE_26_bits),
    .io_connPE_27_ready(continuationNetwork_io_connPE_27_ready),
    .io_connPE_27_valid(continuationNetwork_io_connPE_27_valid),
    .io_connPE_27_bits(continuationNetwork_io_connPE_27_bits),
    .io_connPE_28_ready(continuationNetwork_io_connPE_28_ready),
    .io_connPE_28_valid(continuationNetwork_io_connPE_28_valid),
    .io_connPE_28_bits(continuationNetwork_io_connPE_28_bits),
    .io_connPE_29_ready(continuationNetwork_io_connPE_29_ready),
    .io_connPE_29_valid(continuationNetwork_io_connPE_29_valid),
    .io_connPE_29_bits(continuationNetwork_io_connPE_29_bits),
    .io_connPE_30_ready(continuationNetwork_io_connPE_30_ready),
    .io_connPE_30_valid(continuationNetwork_io_connPE_30_valid),
    .io_connPE_30_bits(continuationNetwork_io_connPE_30_bits),
    .io_connPE_31_ready(continuationNetwork_io_connPE_31_ready),
    .io_connPE_31_valid(continuationNetwork_io_connPE_31_valid),
    .io_connPE_31_bits(continuationNetwork_io_connPE_31_bits),
    .io_connPE_32_ready(continuationNetwork_io_connPE_32_ready),
    .io_connPE_32_valid(continuationNetwork_io_connPE_32_valid),
    .io_connPE_32_bits(continuationNetwork_io_connPE_32_bits),
    .io_connPE_33_ready(continuationNetwork_io_connPE_33_ready),
    .io_connPE_33_valid(continuationNetwork_io_connPE_33_valid),
    .io_connPE_33_bits(continuationNetwork_io_connPE_33_bits),
    .io_connPE_34_ready(continuationNetwork_io_connPE_34_ready),
    .io_connPE_34_valid(continuationNetwork_io_connPE_34_valid),
    .io_connPE_34_bits(continuationNetwork_io_connPE_34_bits),
    .io_connPE_35_ready(continuationNetwork_io_connPE_35_ready),
    .io_connPE_35_valid(continuationNetwork_io_connPE_35_valid),
    .io_connPE_35_bits(continuationNetwork_io_connPE_35_bits),
    .io_connPE_36_ready(continuationNetwork_io_connPE_36_ready),
    .io_connPE_36_valid(continuationNetwork_io_connPE_36_valid),
    .io_connPE_36_bits(continuationNetwork_io_connPE_36_bits),
    .io_connPE_37_ready(continuationNetwork_io_connPE_37_ready),
    .io_connPE_37_valid(continuationNetwork_io_connPE_37_valid),
    .io_connPE_37_bits(continuationNetwork_io_connPE_37_bits),
    .io_connPE_38_ready(continuationNetwork_io_connPE_38_ready),
    .io_connPE_38_valid(continuationNetwork_io_connPE_38_valid),
    .io_connPE_38_bits(continuationNetwork_io_connPE_38_bits),
    .io_connPE_39_ready(continuationNetwork_io_connPE_39_ready),
    .io_connPE_39_valid(continuationNetwork_io_connPE_39_valid),
    .io_connPE_39_bits(continuationNetwork_io_connPE_39_bits),
    .io_connPE_40_ready(continuationNetwork_io_connPE_40_ready),
    .io_connPE_40_valid(continuationNetwork_io_connPE_40_valid),
    .io_connPE_40_bits(continuationNetwork_io_connPE_40_bits),
    .io_connPE_41_ready(continuationNetwork_io_connPE_41_ready),
    .io_connPE_41_valid(continuationNetwork_io_connPE_41_valid),
    .io_connPE_41_bits(continuationNetwork_io_connPE_41_bits),
    .io_connPE_42_ready(continuationNetwork_io_connPE_42_ready),
    .io_connPE_42_valid(continuationNetwork_io_connPE_42_valid),
    .io_connPE_42_bits(continuationNetwork_io_connPE_42_bits),
    .io_connPE_43_ready(continuationNetwork_io_connPE_43_ready),
    .io_connPE_43_valid(continuationNetwork_io_connPE_43_valid),
    .io_connPE_43_bits(continuationNetwork_io_connPE_43_bits),
    .io_connPE_44_ready(continuationNetwork_io_connPE_44_ready),
    .io_connPE_44_valid(continuationNetwork_io_connPE_44_valid),
    .io_connPE_44_bits(continuationNetwork_io_connPE_44_bits),
    .io_connPE_45_ready(continuationNetwork_io_connPE_45_ready),
    .io_connPE_45_valid(continuationNetwork_io_connPE_45_valid),
    .io_connPE_45_bits(continuationNetwork_io_connPE_45_bits),
    .io_connPE_46_ready(continuationNetwork_io_connPE_46_ready),
    .io_connPE_46_valid(continuationNetwork_io_connPE_46_valid),
    .io_connPE_46_bits(continuationNetwork_io_connPE_46_bits),
    .io_connPE_47_ready(continuationNetwork_io_connPE_47_ready),
    .io_connPE_47_valid(continuationNetwork_io_connPE_47_valid),
    .io_connPE_47_bits(continuationNetwork_io_connPE_47_bits),
    .io_connPE_48_ready(continuationNetwork_io_connPE_48_ready),
    .io_connPE_48_valid(continuationNetwork_io_connPE_48_valid),
    .io_connPE_48_bits(continuationNetwork_io_connPE_48_bits),
    .io_connPE_49_ready(continuationNetwork_io_connPE_49_ready),
    .io_connPE_49_valid(continuationNetwork_io_connPE_49_valid),
    .io_connPE_49_bits(continuationNetwork_io_connPE_49_bits),
    .io_connPE_50_ready(continuationNetwork_io_connPE_50_ready),
    .io_connPE_50_valid(continuationNetwork_io_connPE_50_valid),
    .io_connPE_50_bits(continuationNetwork_io_connPE_50_bits),
    .io_connPE_51_ready(continuationNetwork_io_connPE_51_ready),
    .io_connPE_51_valid(continuationNetwork_io_connPE_51_valid),
    .io_connPE_51_bits(continuationNetwork_io_connPE_51_bits),
    .io_connPE_52_ready(continuationNetwork_io_connPE_52_ready),
    .io_connPE_52_valid(continuationNetwork_io_connPE_52_valid),
    .io_connPE_52_bits(continuationNetwork_io_connPE_52_bits),
    .io_connPE_53_ready(continuationNetwork_io_connPE_53_ready),
    .io_connPE_53_valid(continuationNetwork_io_connPE_53_valid),
    .io_connPE_53_bits(continuationNetwork_io_connPE_53_bits),
    .io_connPE_54_ready(continuationNetwork_io_connPE_54_ready),
    .io_connPE_54_valid(continuationNetwork_io_connPE_54_valid),
    .io_connPE_54_bits(continuationNetwork_io_connPE_54_bits),
    .io_connPE_55_ready(continuationNetwork_io_connPE_55_ready),
    .io_connPE_55_valid(continuationNetwork_io_connPE_55_valid),
    .io_connPE_55_bits(continuationNetwork_io_connPE_55_bits),
    .io_connPE_56_ready(continuationNetwork_io_connPE_56_ready),
    .io_connPE_56_valid(continuationNetwork_io_connPE_56_valid),
    .io_connPE_56_bits(continuationNetwork_io_connPE_56_bits),
    .io_connPE_57_ready(continuationNetwork_io_connPE_57_ready),
    .io_connPE_57_valid(continuationNetwork_io_connPE_57_valid),
    .io_connPE_57_bits(continuationNetwork_io_connPE_57_bits),
    .io_connPE_58_ready(continuationNetwork_io_connPE_58_ready),
    .io_connPE_58_valid(continuationNetwork_io_connPE_58_valid),
    .io_connPE_58_bits(continuationNetwork_io_connPE_58_bits),
    .io_connPE_59_ready(continuationNetwork_io_connPE_59_ready),
    .io_connPE_59_valid(continuationNetwork_io_connPE_59_valid),
    .io_connPE_59_bits(continuationNetwork_io_connPE_59_bits),
    .io_connPE_60_ready(continuationNetwork_io_connPE_60_ready),
    .io_connPE_60_valid(continuationNetwork_io_connPE_60_valid),
    .io_connPE_60_bits(continuationNetwork_io_connPE_60_bits),
    .io_connPE_61_ready(continuationNetwork_io_connPE_61_ready),
    .io_connPE_61_valid(continuationNetwork_io_connPE_61_valid),
    .io_connPE_61_bits(continuationNetwork_io_connPE_61_bits),
    .io_connPE_62_ready(continuationNetwork_io_connPE_62_ready),
    .io_connPE_62_valid(continuationNetwork_io_connPE_62_valid),
    .io_connPE_62_bits(continuationNetwork_io_connPE_62_bits),
    .io_connPE_63_ready(continuationNetwork_io_connPE_63_ready),
    .io_connPE_63_valid(continuationNetwork_io_connPE_63_valid),
    .io_connPE_63_bits(continuationNetwork_io_connPE_63_bits)
  );
  virtContAddrServer vcas_0 ( // @[continuationAllocationSide.scala 58:42]
    .clock(vcas_0_clock),
    .reset(vcas_0_reset),
    .io_dataOut_ready(vcas_0_io_dataOut_ready),
    .io_dataOut_valid(vcas_0_io_dataOut_valid),
    .io_dataOut_bits(vcas_0_io_dataOut_bits),
    .io_axi_mgmt_ARREADY(vcas_0_io_axi_mgmt_ARREADY),
    .io_axi_mgmt_ARVALID(vcas_0_io_axi_mgmt_ARVALID),
    .io_axi_mgmt_ARADDR(vcas_0_io_axi_mgmt_ARADDR),
    .io_axi_mgmt_RREADY(vcas_0_io_axi_mgmt_RREADY),
    .io_axi_mgmt_RVALID(vcas_0_io_axi_mgmt_RVALID),
    .io_axi_mgmt_RDATA(vcas_0_io_axi_mgmt_RDATA),
    .io_axi_mgmt_AWREADY(vcas_0_io_axi_mgmt_AWREADY),
    .io_axi_mgmt_AWVALID(vcas_0_io_axi_mgmt_AWVALID),
    .io_axi_mgmt_AWADDR(vcas_0_io_axi_mgmt_AWADDR),
    .io_axi_mgmt_WREADY(vcas_0_io_axi_mgmt_WREADY),
    .io_axi_mgmt_WVALID(vcas_0_io_axi_mgmt_WVALID),
    .io_axi_mgmt_WDATA(vcas_0_io_axi_mgmt_WDATA),
    .io_axi_mgmt_WSTRB(vcas_0_io_axi_mgmt_WSTRB),
    .io_axi_mgmt_BREADY(vcas_0_io_axi_mgmt_BREADY),
    .io_axi_mgmt_BVALID(vcas_0_io_axi_mgmt_BVALID),
    .io_read_address_ready(vcas_0_io_read_address_ready),
    .io_read_address_valid(vcas_0_io_read_address_valid),
    .io_read_address_bits(vcas_0_io_read_address_bits),
    .io_read_data_ready(vcas_0_io_read_data_ready),
    .io_read_data_valid(vcas_0_io_read_data_valid),
    .io_read_data_bits(vcas_0_io_read_data_bits)
  );
  readyValidMem_1 vcasRvmRO_0 ( // @[continuationAllocationSide.scala 71:47]
    .io_read_address_ready(vcasRvmRO_0_io_read_address_ready),
    .io_read_address_valid(vcasRvmRO_0_io_read_address_valid),
    .io_read_address_bits(vcasRvmRO_0_io_read_address_bits),
    .io_read_data_ready(vcasRvmRO_0_io_read_data_ready),
    .io_read_data_valid(vcasRvmRO_0_io_read_data_valid),
    .io_read_data_bits(vcasRvmRO_0_io_read_data_bits),
    .axi_ARREADY(vcasRvmRO_0_axi_ARREADY),
    .axi_ARVALID(vcasRvmRO_0_axi_ARVALID),
    .axi_ARADDR(vcasRvmRO_0_axi_ARADDR),
    .axi_RREADY(vcasRvmRO_0_axi_RREADY),
    .axi_RVALID(vcasRvmRO_0_axi_RVALID),
    .axi_RDATA(vcasRvmRO_0_axi_RDATA)
  );
  assign io_contOut_0_TVALID = continuationNetwork_io_connPE_0_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_0_TDATA = continuationNetwork_io_connPE_0_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_1_TVALID = continuationNetwork_io_connPE_1_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_1_TDATA = continuationNetwork_io_connPE_1_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_2_TVALID = continuationNetwork_io_connPE_2_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_2_TDATA = continuationNetwork_io_connPE_2_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_3_TVALID = continuationNetwork_io_connPE_3_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_3_TDATA = continuationNetwork_io_connPE_3_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_4_TVALID = continuationNetwork_io_connPE_4_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_4_TDATA = continuationNetwork_io_connPE_4_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_5_TVALID = continuationNetwork_io_connPE_5_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_5_TDATA = continuationNetwork_io_connPE_5_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_6_TVALID = continuationNetwork_io_connPE_6_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_6_TDATA = continuationNetwork_io_connPE_6_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_7_TVALID = continuationNetwork_io_connPE_7_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_7_TDATA = continuationNetwork_io_connPE_7_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_8_TVALID = continuationNetwork_io_connPE_8_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_8_TDATA = continuationNetwork_io_connPE_8_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_9_TVALID = continuationNetwork_io_connPE_9_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_9_TDATA = continuationNetwork_io_connPE_9_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_10_TVALID = continuationNetwork_io_connPE_10_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_10_TDATA = continuationNetwork_io_connPE_10_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_11_TVALID = continuationNetwork_io_connPE_11_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_11_TDATA = continuationNetwork_io_connPE_11_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_12_TVALID = continuationNetwork_io_connPE_12_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_12_TDATA = continuationNetwork_io_connPE_12_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_13_TVALID = continuationNetwork_io_connPE_13_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_13_TDATA = continuationNetwork_io_connPE_13_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_14_TVALID = continuationNetwork_io_connPE_14_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_14_TDATA = continuationNetwork_io_connPE_14_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_15_TVALID = continuationNetwork_io_connPE_15_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_15_TDATA = continuationNetwork_io_connPE_15_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_16_TVALID = continuationNetwork_io_connPE_16_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_16_TDATA = continuationNetwork_io_connPE_16_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_17_TVALID = continuationNetwork_io_connPE_17_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_17_TDATA = continuationNetwork_io_connPE_17_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_18_TVALID = continuationNetwork_io_connPE_18_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_18_TDATA = continuationNetwork_io_connPE_18_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_19_TVALID = continuationNetwork_io_connPE_19_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_19_TDATA = continuationNetwork_io_connPE_19_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_20_TVALID = continuationNetwork_io_connPE_20_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_20_TDATA = continuationNetwork_io_connPE_20_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_21_TVALID = continuationNetwork_io_connPE_21_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_21_TDATA = continuationNetwork_io_connPE_21_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_22_TVALID = continuationNetwork_io_connPE_22_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_22_TDATA = continuationNetwork_io_connPE_22_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_23_TVALID = continuationNetwork_io_connPE_23_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_23_TDATA = continuationNetwork_io_connPE_23_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_24_TVALID = continuationNetwork_io_connPE_24_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_24_TDATA = continuationNetwork_io_connPE_24_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_25_TVALID = continuationNetwork_io_connPE_25_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_25_TDATA = continuationNetwork_io_connPE_25_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_26_TVALID = continuationNetwork_io_connPE_26_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_26_TDATA = continuationNetwork_io_connPE_26_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_27_TVALID = continuationNetwork_io_connPE_27_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_27_TDATA = continuationNetwork_io_connPE_27_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_28_TVALID = continuationNetwork_io_connPE_28_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_28_TDATA = continuationNetwork_io_connPE_28_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_29_TVALID = continuationNetwork_io_connPE_29_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_29_TDATA = continuationNetwork_io_connPE_29_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_30_TVALID = continuationNetwork_io_connPE_30_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_30_TDATA = continuationNetwork_io_connPE_30_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_31_TVALID = continuationNetwork_io_connPE_31_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_31_TDATA = continuationNetwork_io_connPE_31_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_32_TVALID = continuationNetwork_io_connPE_32_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_32_TDATA = continuationNetwork_io_connPE_32_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_33_TVALID = continuationNetwork_io_connPE_33_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_33_TDATA = continuationNetwork_io_connPE_33_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_34_TVALID = continuationNetwork_io_connPE_34_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_34_TDATA = continuationNetwork_io_connPE_34_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_35_TVALID = continuationNetwork_io_connPE_35_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_35_TDATA = continuationNetwork_io_connPE_35_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_36_TVALID = continuationNetwork_io_connPE_36_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_36_TDATA = continuationNetwork_io_connPE_36_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_37_TVALID = continuationNetwork_io_connPE_37_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_37_TDATA = continuationNetwork_io_connPE_37_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_38_TVALID = continuationNetwork_io_connPE_38_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_38_TDATA = continuationNetwork_io_connPE_38_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_39_TVALID = continuationNetwork_io_connPE_39_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_39_TDATA = continuationNetwork_io_connPE_39_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_40_TVALID = continuationNetwork_io_connPE_40_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_40_TDATA = continuationNetwork_io_connPE_40_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_41_TVALID = continuationNetwork_io_connPE_41_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_41_TDATA = continuationNetwork_io_connPE_41_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_42_TVALID = continuationNetwork_io_connPE_42_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_42_TDATA = continuationNetwork_io_connPE_42_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_43_TVALID = continuationNetwork_io_connPE_43_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_43_TDATA = continuationNetwork_io_connPE_43_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_44_TVALID = continuationNetwork_io_connPE_44_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_44_TDATA = continuationNetwork_io_connPE_44_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_45_TVALID = continuationNetwork_io_connPE_45_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_45_TDATA = continuationNetwork_io_connPE_45_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_46_TVALID = continuationNetwork_io_connPE_46_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_46_TDATA = continuationNetwork_io_connPE_46_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_47_TVALID = continuationNetwork_io_connPE_47_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_47_TDATA = continuationNetwork_io_connPE_47_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_48_TVALID = continuationNetwork_io_connPE_48_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_48_TDATA = continuationNetwork_io_connPE_48_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_49_TVALID = continuationNetwork_io_connPE_49_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_49_TDATA = continuationNetwork_io_connPE_49_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_50_TVALID = continuationNetwork_io_connPE_50_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_50_TDATA = continuationNetwork_io_connPE_50_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_51_TVALID = continuationNetwork_io_connPE_51_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_51_TDATA = continuationNetwork_io_connPE_51_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_52_TVALID = continuationNetwork_io_connPE_52_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_52_TDATA = continuationNetwork_io_connPE_52_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_53_TVALID = continuationNetwork_io_connPE_53_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_53_TDATA = continuationNetwork_io_connPE_53_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_54_TVALID = continuationNetwork_io_connPE_54_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_54_TDATA = continuationNetwork_io_connPE_54_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_55_TVALID = continuationNetwork_io_connPE_55_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_55_TDATA = continuationNetwork_io_connPE_55_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_56_TVALID = continuationNetwork_io_connPE_56_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_56_TDATA = continuationNetwork_io_connPE_56_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_57_TVALID = continuationNetwork_io_connPE_57_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_57_TDATA = continuationNetwork_io_connPE_57_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_58_TVALID = continuationNetwork_io_connPE_58_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_58_TDATA = continuationNetwork_io_connPE_58_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_59_TVALID = continuationNetwork_io_connPE_59_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_59_TDATA = continuationNetwork_io_connPE_59_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_60_TVALID = continuationNetwork_io_connPE_60_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_60_TDATA = continuationNetwork_io_connPE_60_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_61_TVALID = continuationNetwork_io_connPE_61_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_61_TDATA = continuationNetwork_io_connPE_61_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_62_TVALID = continuationNetwork_io_connPE_62_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_62_TDATA = continuationNetwork_io_connPE_62_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_63_TVALID = continuationNetwork_io_connPE_63_valid; // @[continuationAllocationSide.scala 85:42]
  assign io_contOut_63_TDATA = continuationNetwork_io_connPE_63_bits; // @[continuationAllocationSide.scala 85:42]
  assign io_axi_mgmt_vcas_0_ARREADY = vcas_0_io_axi_mgmt_ARREADY; // @[continuationAllocationSide.scala 75:43]
  assign io_axi_mgmt_vcas_0_RVALID = vcas_0_io_axi_mgmt_RVALID; // @[continuationAllocationSide.scala 75:43]
  assign io_axi_mgmt_vcas_0_RDATA = vcas_0_io_axi_mgmt_RDATA; // @[continuationAllocationSide.scala 75:43]
  assign io_axi_mgmt_vcas_0_AWREADY = vcas_0_io_axi_mgmt_AWREADY; // @[continuationAllocationSide.scala 75:43]
  assign io_axi_mgmt_vcas_0_WREADY = vcas_0_io_axi_mgmt_WREADY; // @[continuationAllocationSide.scala 75:43]
  assign io_axi_mgmt_vcas_0_BVALID = vcas_0_io_axi_mgmt_BVALID; // @[continuationAllocationSide.scala 75:43]
  assign io_vcas_axi_full_0_ARVALID = vcasRvmRO_0_axi_ARVALID; // @[continuationAllocationSide.scala 79:43]
  assign io_vcas_axi_full_0_ARADDR = vcasRvmRO_0_axi_ARADDR; // @[continuationAllocationSide.scala 79:43]
  assign io_vcas_axi_full_0_RREADY = vcasRvmRO_0_axi_RREADY; // @[continuationAllocationSide.scala 79:43]
  assign continuationNetwork_clock = clock;
  assign continuationNetwork_reset = reset;
  assign continuationNetwork_io_connVCAS_0_valid = vcas_0_io_dataOut_valid; // @[continuationAllocationSide.scala 80:45]
  assign continuationNetwork_io_connVCAS_0_bits = vcas_0_io_dataOut_bits; // @[continuationAllocationSide.scala 80:45]
  assign continuationNetwork_io_connPE_0_ready = io_contOut_0_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_1_ready = io_contOut_1_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_2_ready = io_contOut_2_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_3_ready = io_contOut_3_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_4_ready = io_contOut_4_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_5_ready = io_contOut_5_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_6_ready = io_contOut_6_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_7_ready = io_contOut_7_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_8_ready = io_contOut_8_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_9_ready = io_contOut_9_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_10_ready = io_contOut_10_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_11_ready = io_contOut_11_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_12_ready = io_contOut_12_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_13_ready = io_contOut_13_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_14_ready = io_contOut_14_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_15_ready = io_contOut_15_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_16_ready = io_contOut_16_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_17_ready = io_contOut_17_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_18_ready = io_contOut_18_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_19_ready = io_contOut_19_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_20_ready = io_contOut_20_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_21_ready = io_contOut_21_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_22_ready = io_contOut_22_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_23_ready = io_contOut_23_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_24_ready = io_contOut_24_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_25_ready = io_contOut_25_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_26_ready = io_contOut_26_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_27_ready = io_contOut_27_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_28_ready = io_contOut_28_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_29_ready = io_contOut_29_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_30_ready = io_contOut_30_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_31_ready = io_contOut_31_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_32_ready = io_contOut_32_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_33_ready = io_contOut_33_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_34_ready = io_contOut_34_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_35_ready = io_contOut_35_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_36_ready = io_contOut_36_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_37_ready = io_contOut_37_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_38_ready = io_contOut_38_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_39_ready = io_contOut_39_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_40_ready = io_contOut_40_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_41_ready = io_contOut_41_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_42_ready = io_contOut_42_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_43_ready = io_contOut_43_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_44_ready = io_contOut_44_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_45_ready = io_contOut_45_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_46_ready = io_contOut_46_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_47_ready = io_contOut_47_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_48_ready = io_contOut_48_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_49_ready = io_contOut_49_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_50_ready = io_contOut_50_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_51_ready = io_contOut_51_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_52_ready = io_contOut_52_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_53_ready = io_contOut_53_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_54_ready = io_contOut_54_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_55_ready = io_contOut_55_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_56_ready = io_contOut_56_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_57_ready = io_contOut_57_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_58_ready = io_contOut_58_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_59_ready = io_contOut_59_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_60_ready = io_contOut_60_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_61_ready = io_contOut_61_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_62_ready = io_contOut_62_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign continuationNetwork_io_connPE_63_ready = io_contOut_63_TREADY; // @[continuationAllocationSide.scala 85:42]
  assign vcas_0_clock = clock;
  assign vcas_0_reset = reset;
  assign vcas_0_io_dataOut_ready = continuationNetwork_io_connVCAS_0_ready; // @[continuationAllocationSide.scala 80:45]
  assign vcas_0_io_axi_mgmt_ARVALID = io_axi_mgmt_vcas_0_ARVALID; // @[continuationAllocationSide.scala 75:43]
  assign vcas_0_io_axi_mgmt_ARADDR = io_axi_mgmt_vcas_0_ARADDR; // @[continuationAllocationSide.scala 75:43]
  assign vcas_0_io_axi_mgmt_RREADY = io_axi_mgmt_vcas_0_RREADY; // @[continuationAllocationSide.scala 75:43]
  assign vcas_0_io_axi_mgmt_AWVALID = io_axi_mgmt_vcas_0_AWVALID; // @[continuationAllocationSide.scala 75:43]
  assign vcas_0_io_axi_mgmt_AWADDR = io_axi_mgmt_vcas_0_AWADDR; // @[continuationAllocationSide.scala 75:43]
  assign vcas_0_io_axi_mgmt_WVALID = io_axi_mgmt_vcas_0_WVALID; // @[continuationAllocationSide.scala 75:43]
  assign vcas_0_io_axi_mgmt_WDATA = io_axi_mgmt_vcas_0_WDATA; // @[continuationAllocationSide.scala 75:43]
  assign vcas_0_io_axi_mgmt_WSTRB = io_axi_mgmt_vcas_0_WSTRB; // @[continuationAllocationSide.scala 75:43]
  assign vcas_0_io_axi_mgmt_BREADY = io_axi_mgmt_vcas_0_BREADY; // @[continuationAllocationSide.scala 75:43]
  assign vcas_0_io_read_address_ready = vcasRvmRO_0_io_read_address_ready; // @[continuationAllocationSide.scala 77:43]
  assign vcas_0_io_read_data_valid = vcasRvmRO_0_io_read_data_valid; // @[continuationAllocationSide.scala 78:43]
  assign vcas_0_io_read_data_bits = vcasRvmRO_0_io_read_data_bits; // @[continuationAllocationSide.scala 78:43]
  assign vcasRvmRO_0_io_read_address_valid = vcas_0_io_read_address_valid; // @[continuationAllocationSide.scala 77:43]
  assign vcasRvmRO_0_io_read_address_bits = vcas_0_io_read_address_bits; // @[continuationAllocationSide.scala 77:43]
  assign vcasRvmRO_0_io_read_data_ready = vcas_0_io_read_data_ready; // @[continuationAllocationSide.scala 78:43]
  assign vcasRvmRO_0_axi_ARREADY = io_vcas_axi_full_0_ARREADY; // @[continuationAllocationSide.scala 79:43]
  assign vcasRvmRO_0_axi_RVALID = io_vcas_axi_full_0_RVALID; // @[continuationAllocationSide.scala 79:43]
  assign vcasRvmRO_0_axi_RDATA = io_vcas_axi_full_0_RDATA; // @[continuationAllocationSide.scala 79:43]
endmodule
module argRouteNtwUnit(
  input         clock,
  input         reset,
  output        io_addressIn_ready,
  input         io_addressIn_valid,
  input  [63:0] io_addressIn_bits,
  output        io_peAddress_ready,
  input         io_peAddress_valid,
  input  [63:0] io_peAddress_bits,
  input         io_addressOut_ready,
  output        io_addressOut_valid,
  output [63:0] io_addressOut_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  stateReg; // @[argRouteNtwUnit.scala 22:30]
  reg [63:0] addressReg; // @[argRouteNtwUnit.scala 23:30]
  reg  priorityReg; // @[argRouteNtwUnit.scala 24:30]
  wire  _T = ~stateReg; // @[argRouteNtwUnit.scala 33:19]
  wire  _T_1 = io_addressIn_valid & io_peAddress_valid; // @[argRouteNtwUnit.scala 34:33]
  wire [63:0] _GEN_1 = io_addressIn_valid ? io_addressIn_bits : addressReg; // @[argRouteNtwUnit.scala 44:43 45:28 23:30]
  wire  _GEN_4 = io_addressIn_valid & io_peAddress_valid ? ~priorityReg : priorityReg; // @[argRouteNtwUnit.scala 34:55 40:25 24:30]
  wire  _GEN_5 = io_addressIn_valid | io_peAddress_valid | stateReg; // @[argRouteNtwUnit.scala 49:55 50:24 22:30]
  wire  _GEN_6 = io_addressOut_ready ? 1'h0 : stateReg; // @[argRouteNtwUnit.scala 54:34 55:22 22:30]
  wire  _GEN_7 = stateReg & _GEN_6; // @[argRouteNtwUnit.scala 53:44 58:18]
  wire  _GEN_9 = ~stateReg ? _GEN_4 : priorityReg; // @[argRouteNtwUnit.scala 24:30 33:43]
  wire  _GEN_12 = priorityReg ? 1'h0 : 1'h1; // @[argRouteNtwUnit.scala 26:28 64:30 67:36]
  wire  _GEN_15 = io_peAddress_valid ? 1'h0 : io_addressIn_valid; // @[argRouteNtwUnit.scala 26:28 70:37]
  wire  _GEN_16 = _T_1 ? priorityReg : io_peAddress_valid; // @[argRouteNtwUnit.scala 63:55]
  wire  _GEN_17 = _T_1 ? _GEN_12 : _GEN_15; // @[argRouteNtwUnit.scala 63:55]
  assign io_addressIn_ready = _T & _GEN_17; // @[argRouteNtwUnit.scala 26:28 62:43]
  assign io_peAddress_ready = _T & _GEN_16; // @[argRouteNtwUnit.scala 27:28 62:43]
  assign io_addressOut_valid = _T ? 1'h0 : stateReg; // @[argRouteNtwUnit.scala 28:28 62:43]
  assign io_addressOut_bits = addressReg; // @[argRouteNtwUnit.scala 29:28]
  always @(posedge clock) begin
    if (reset) begin // @[argRouteNtwUnit.scala 22:30]
      stateReg <= 1'h0; // @[argRouteNtwUnit.scala 22:30]
    end else if (~stateReg) begin // @[argRouteNtwUnit.scala 33:43]
      stateReg <= _GEN_5;
    end else begin
      stateReg <= _GEN_7;
    end
    if (reset) begin // @[argRouteNtwUnit.scala 23:30]
      addressReg <= 64'h0; // @[argRouteNtwUnit.scala 23:30]
    end else if (~stateReg) begin // @[argRouteNtwUnit.scala 33:43]
      if (io_addressIn_valid & io_peAddress_valid) begin // @[argRouteNtwUnit.scala 34:55]
        if (priorityReg) begin // @[argRouteNtwUnit.scala 35:30]
          addressReg <= io_peAddress_bits; // @[argRouteNtwUnit.scala 36:28]
        end else begin
          addressReg <= io_addressIn_bits; // @[argRouteNtwUnit.scala 38:28]
        end
      end else if (io_peAddress_valid) begin // @[argRouteNtwUnit.scala 42:37]
        addressReg <= io_peAddress_bits; // @[argRouteNtwUnit.scala 43:28]
      end else begin
        addressReg <= _GEN_1;
      end
    end
    priorityReg <= reset | _GEN_9; // @[argRouteNtwUnit.scala 24:{30,30}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  addressReg = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  priorityReg = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module argRouteNtwVirtUnit(
  input         clock,
  input         reset,
  output        io_addressIn_ready,
  input         io_addressIn_valid,
  input  [63:0] io_addressIn_bits,
  input         io_vasAddressOut_ready,
  output        io_vasAddressOut_valid,
  output [63:0] io_vasAddressOut_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] stateReg; // @[argRouteNtwVirtUnit.scala 23:32]
  reg [63:0] addressReg; // @[argRouteNtwVirtUnit.scala 24:32]
  wire [1:0] mask = 2'h2 - 2'h1; // @[argRouteNtwVirtUnit.scala 25:49]
  wire  _T = stateReg == 2'h0; // @[argRouteNtwVirtUnit.scala 33:19]
  wire [58:0] _GEN_7 = {{57'd0}, mask}; // @[argRouteNtwVirtUnit.scala 45:57]
  wire [58:0] _T_2 = io_addressIn_bits[63:5] & _GEN_7; // @[argRouteNtwVirtUnit.scala 45:57]
  wire  _T_4 = stateReg == 2'h1; // @[argRouteNtwVirtUnit.scala 52:25]
  wire  _T_5 = stateReg == 2'h2; // @[argRouteNtwVirtUnit.scala 57:25]
  wire [1:0] _GEN_4 = io_vasAddressOut_ready ? 2'h0 : stateReg; // @[argRouteNtwVirtUnit.scala 59:37 60:22 23:32]
  wire  _GEN_9 = stateReg == 2'h1 ? 1'h0 : _T_5; // @[argRouteNtwVirtUnit.scala 28:28 52:48]
  wire  _GEN_14 = stateReg == 2'h0 ? 1'h0 : _GEN_9; // @[argRouteNtwVirtUnit.scala 28:28 33:43]
  wire  _GEN_15 = _T_5 | _GEN_14; // @[argRouteNtwVirtUnit.scala 68:47 69:32]
  wire  _GEN_17 = _T_4 ? _GEN_14 : _GEN_15; // @[argRouteNtwVirtUnit.scala 66:48]
  assign io_addressIn_ready = _T | _T; // @[argRouteNtwVirtUnit.scala 64:43 65:28]
  assign io_vasAddressOut_valid = _T ? _GEN_14 : _GEN_17; // @[argRouteNtwVirtUnit.scala 64:43]
  assign io_vasAddressOut_bits = addressReg; // @[argRouteNtwVirtUnit.scala 30:28]
  always @(posedge clock) begin
    if (reset) begin // @[argRouteNtwVirtUnit.scala 23:32]
      stateReg <= 2'h0; // @[argRouteNtwVirtUnit.scala 23:32]
    end else if (stateReg == 2'h0) begin // @[argRouteNtwVirtUnit.scala 33:43]
      if (io_addressIn_valid) begin // @[argRouteNtwVirtUnit.scala 35:33]
        if (_T_2 == 59'h0) begin // @[argRouteNtwVirtUnit.scala 45:104]
          stateReg <= 2'h2; // @[argRouteNtwVirtUnit.scala 46:30]
        end else begin
          stateReg <= 2'h1; // @[argRouteNtwVirtUnit.scala 48:30]
        end
      end
    end else if (!(stateReg == 2'h1)) begin // @[argRouteNtwVirtUnit.scala 52:48]
      if (stateReg == 2'h2) begin // @[argRouteNtwVirtUnit.scala 57:47]
        stateReg <= _GEN_4;
      end
    end
    if (reset) begin // @[argRouteNtwVirtUnit.scala 24:32]
      addressReg <= 64'h0; // @[argRouteNtwVirtUnit.scala 24:32]
    end else if (stateReg == 2'h0) begin // @[argRouteNtwVirtUnit.scala 33:43]
      if (io_addressIn_valid) begin // @[argRouteNtwVirtUnit.scala 35:33]
        addressReg <= io_addressIn_bits; // @[argRouteNtwVirtUnit.scala 36:24]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  addressReg = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module argRouteNtwVirtUnit_1(
  input         clock,
  input         reset,
  output        io_addressIn_ready,
  input         io_addressIn_valid,
  input  [63:0] io_addressIn_bits,
  input         io_vasAddressOut_ready,
  output        io_vasAddressOut_valid,
  output [63:0] io_vasAddressOut_bits,
  input         io_addressOut_ready,
  output        io_addressOut_valid,
  output [63:0] io_addressOut_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] stateReg; // @[argRouteNtwVirtUnit.scala 23:32]
  reg [63:0] addressReg; // @[argRouteNtwVirtUnit.scala 24:32]
  wire [1:0] mask = 2'h2 - 2'h1; // @[argRouteNtwVirtUnit.scala 25:49]
  wire  _T = stateReg == 2'h0; // @[argRouteNtwVirtUnit.scala 33:19]
  wire [58:0] _GEN_21 = {{57'd0}, mask}; // @[argRouteNtwVirtUnit.scala 45:57]
  wire [58:0] _T_2 = io_addressIn_bits[63:5] & _GEN_21; // @[argRouteNtwVirtUnit.scala 45:57]
  wire  _T_4 = stateReg == 2'h1; // @[argRouteNtwVirtUnit.scala 52:25]
  wire  _T_5 = stateReg == 2'h2; // @[argRouteNtwVirtUnit.scala 57:25]
  wire [1:0] _GEN_4 = io_vasAddressOut_ready ? 2'h0 : stateReg; // @[argRouteNtwVirtUnit.scala 59:37 60:22 23:32]
  wire  _GEN_9 = stateReg == 2'h1 ? 1'h0 : _T_5; // @[argRouteNtwVirtUnit.scala 28:28 52:48]
  wire  _GEN_13 = stateReg == 2'h0 ? 1'h0 : _T_4; // @[argRouteNtwVirtUnit.scala 29:28 33:43]
  wire  _GEN_14 = stateReg == 2'h0 ? 1'h0 : _GEN_9; // @[argRouteNtwVirtUnit.scala 28:28 33:43]
  wire  _GEN_15 = _T_5 | _GEN_14; // @[argRouteNtwVirtUnit.scala 68:47 69:32]
  wire  _GEN_16 = _T_4 | _GEN_13; // @[argRouteNtwVirtUnit.scala 66:48 67:29]
  wire  _GEN_17 = _T_4 ? _GEN_14 : _GEN_15; // @[argRouteNtwVirtUnit.scala 66:48]
  assign io_addressIn_ready = _T | _T; // @[argRouteNtwVirtUnit.scala 64:43 65:28]
  assign io_vasAddressOut_valid = _T ? _GEN_14 : _GEN_17; // @[argRouteNtwVirtUnit.scala 64:43]
  assign io_vasAddressOut_bits = addressReg; // @[argRouteNtwVirtUnit.scala 30:28]
  assign io_addressOut_valid = _T ? _GEN_13 : _GEN_16; // @[argRouteNtwVirtUnit.scala 64:43]
  assign io_addressOut_bits = addressReg; // @[argRouteNtwVirtUnit.scala 31:28]
  always @(posedge clock) begin
    if (reset) begin // @[argRouteNtwVirtUnit.scala 23:32]
      stateReg <= 2'h0; // @[argRouteNtwVirtUnit.scala 23:32]
    end else if (stateReg == 2'h0) begin // @[argRouteNtwVirtUnit.scala 33:43]
      if (io_addressIn_valid) begin // @[argRouteNtwVirtUnit.scala 35:33]
        if (_T_2 == 59'h1) begin // @[argRouteNtwVirtUnit.scala 45:104]
          stateReg <= 2'h2; // @[argRouteNtwVirtUnit.scala 46:30]
        end else begin
          stateReg <= 2'h1; // @[argRouteNtwVirtUnit.scala 48:30]
        end
      end
    end else if (stateReg == 2'h1) begin // @[argRouteNtwVirtUnit.scala 52:48]
      if (io_addressOut_ready) begin // @[argRouteNtwVirtUnit.scala 54:34]
        stateReg <= 2'h0; // @[argRouteNtwVirtUnit.scala 55:22]
      end
    end else if (stateReg == 2'h2) begin // @[argRouteNtwVirtUnit.scala 57:47]
      stateReg <= _GEN_4;
    end
    if (reset) begin // @[argRouteNtwVirtUnit.scala 24:32]
      addressReg <= 64'h0; // @[argRouteNtwVirtUnit.scala 24:32]
    end else if (stateReg == 2'h0) begin // @[argRouteNtwVirtUnit.scala 33:43]
      if (io_addressIn_valid) begin // @[argRouteNtwVirtUnit.scala 35:33]
        addressReg <= io_addressIn_bits; // @[argRouteNtwVirtUnit.scala 36:24]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  addressReg = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_71(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram [0:31]; // @[Decoupled.scala 275:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 275:95]
  wire [4:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 275:95]
  wire [63:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 275:95]
  wire [63:0] ram_MPORT_data; // @[Decoupled.scala 275:95]
  wire [4:0] ram_MPORT_addr; // @[Decoupled.scala 275:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 275:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 275:95]
  reg [4:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [4:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 278:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 279:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 280:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 281:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 52:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 52:35]
  wire [4:0] _value_T_1 = enq_ptr_value + 5'h1; // @[Counter.scala 77:24]
  wire [4:0] _value_T_3 = deq_ptr_value + 5'h1; // @[Counter.scala 77:24]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 275:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 305:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 304:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 312:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 275:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 5'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 288:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 5'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 292:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 278:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 278:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 295:27]
      maybe_full <= do_enq; // @[Decoupled.scala 296:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module contQueue_64(
  input         clock,
  input         reset,
  output        io_addressIn_ready,
  input         io_addressIn_valid,
  input  [63:0] io_addressIn_bits,
  input         io_addressOut_ready,
  output        io_addressOut_valid,
  output [63:0] io_addressOut_bits
);
  wire  q_clock; // @[contQueue.scala 13:19]
  wire  q_reset; // @[contQueue.scala 13:19]
  wire  q_io_enq_ready; // @[contQueue.scala 13:19]
  wire  q_io_enq_valid; // @[contQueue.scala 13:19]
  wire [63:0] q_io_enq_bits; // @[contQueue.scala 13:19]
  wire  q_io_deq_ready; // @[contQueue.scala 13:19]
  wire  q_io_deq_valid; // @[contQueue.scala 13:19]
  wire [63:0] q_io_deq_bits; // @[contQueue.scala 13:19]
  Queue_71 q ( // @[contQueue.scala 13:19]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits(q_io_enq_bits),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits(q_io_deq_bits)
  );
  assign io_addressIn_ready = q_io_enq_ready; // @[contQueue.scala 15:14]
  assign io_addressOut_valid = q_io_deq_valid; // @[contQueue.scala 16:19]
  assign io_addressOut_bits = q_io_deq_bits; // @[contQueue.scala 16:19]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_addressIn_valid; // @[contQueue.scala 15:14]
  assign q_io_enq_bits = io_addressIn_bits; // @[contQueue.scala 15:14]
  assign q_io_deq_ready = io_addressOut_ready; // @[contQueue.scala 16:19]
endmodule
module argRouteNetwork(
  input         clock,
  input         reset,
  input         io_connVAS_0_ready,
  output        io_connVAS_0_valid,
  output [63:0] io_connVAS_0_bits,
  input         io_connVAS_1_ready,
  output        io_connVAS_1_valid,
  output [63:0] io_connVAS_1_bits,
  output        io_connPE_0_ready,
  input         io_connPE_0_valid,
  input  [63:0] io_connPE_0_bits,
  output        io_connPE_1_ready,
  input         io_connPE_1_valid,
  input  [63:0] io_connPE_1_bits,
  output        io_connPE_2_ready,
  input         io_connPE_2_valid,
  input  [63:0] io_connPE_2_bits,
  output        io_connPE_3_ready,
  input         io_connPE_3_valid,
  input  [63:0] io_connPE_3_bits,
  output        io_connPE_4_ready,
  input         io_connPE_4_valid,
  input  [63:0] io_connPE_4_bits,
  output        io_connPE_5_ready,
  input         io_connPE_5_valid,
  input  [63:0] io_connPE_5_bits,
  output        io_connPE_6_ready,
  input         io_connPE_6_valid,
  input  [63:0] io_connPE_6_bits,
  output        io_connPE_7_ready,
  input         io_connPE_7_valid,
  input  [63:0] io_connPE_7_bits,
  output        io_connPE_8_ready,
  input         io_connPE_8_valid,
  input  [63:0] io_connPE_8_bits,
  output        io_connPE_9_ready,
  input         io_connPE_9_valid,
  input  [63:0] io_connPE_9_bits,
  output        io_connPE_10_ready,
  input         io_connPE_10_valid,
  input  [63:0] io_connPE_10_bits,
  output        io_connPE_11_ready,
  input         io_connPE_11_valid,
  input  [63:0] io_connPE_11_bits,
  output        io_connPE_12_ready,
  input         io_connPE_12_valid,
  input  [63:0] io_connPE_12_bits,
  output        io_connPE_13_ready,
  input         io_connPE_13_valid,
  input  [63:0] io_connPE_13_bits,
  output        io_connPE_14_ready,
  input         io_connPE_14_valid,
  input  [63:0] io_connPE_14_bits,
  output        io_connPE_15_ready,
  input         io_connPE_15_valid,
  input  [63:0] io_connPE_15_bits,
  output        io_connPE_16_ready,
  input         io_connPE_16_valid,
  input  [63:0] io_connPE_16_bits,
  output        io_connPE_17_ready,
  input         io_connPE_17_valid,
  input  [63:0] io_connPE_17_bits,
  output        io_connPE_18_ready,
  input         io_connPE_18_valid,
  input  [63:0] io_connPE_18_bits,
  output        io_connPE_19_ready,
  input         io_connPE_19_valid,
  input  [63:0] io_connPE_19_bits,
  output        io_connPE_20_ready,
  input         io_connPE_20_valid,
  input  [63:0] io_connPE_20_bits,
  output        io_connPE_21_ready,
  input         io_connPE_21_valid,
  input  [63:0] io_connPE_21_bits,
  output        io_connPE_22_ready,
  input         io_connPE_22_valid,
  input  [63:0] io_connPE_22_bits,
  output        io_connPE_23_ready,
  input         io_connPE_23_valid,
  input  [63:0] io_connPE_23_bits,
  output        io_connPE_24_ready,
  input         io_connPE_24_valid,
  input  [63:0] io_connPE_24_bits,
  output        io_connPE_25_ready,
  input         io_connPE_25_valid,
  input  [63:0] io_connPE_25_bits,
  output        io_connPE_26_ready,
  input         io_connPE_26_valid,
  input  [63:0] io_connPE_26_bits,
  output        io_connPE_27_ready,
  input         io_connPE_27_valid,
  input  [63:0] io_connPE_27_bits,
  output        io_connPE_28_ready,
  input         io_connPE_28_valid,
  input  [63:0] io_connPE_28_bits,
  output        io_connPE_29_ready,
  input         io_connPE_29_valid,
  input  [63:0] io_connPE_29_bits,
  output        io_connPE_30_ready,
  input         io_connPE_30_valid,
  input  [63:0] io_connPE_30_bits,
  output        io_connPE_31_ready,
  input         io_connPE_31_valid,
  input  [63:0] io_connPE_31_bits,
  output        io_connPE_32_ready,
  input         io_connPE_32_valid,
  input  [63:0] io_connPE_32_bits,
  output        io_connPE_33_ready,
  input         io_connPE_33_valid,
  input  [63:0] io_connPE_33_bits,
  output        io_connPE_34_ready,
  input         io_connPE_34_valid,
  input  [63:0] io_connPE_34_bits,
  output        io_connPE_35_ready,
  input         io_connPE_35_valid,
  input  [63:0] io_connPE_35_bits,
  output        io_connPE_36_ready,
  input         io_connPE_36_valid,
  input  [63:0] io_connPE_36_bits,
  output        io_connPE_37_ready,
  input         io_connPE_37_valid,
  input  [63:0] io_connPE_37_bits,
  output        io_connPE_38_ready,
  input         io_connPE_38_valid,
  input  [63:0] io_connPE_38_bits,
  output        io_connPE_39_ready,
  input         io_connPE_39_valid,
  input  [63:0] io_connPE_39_bits,
  output        io_connPE_40_ready,
  input         io_connPE_40_valid,
  input  [63:0] io_connPE_40_bits,
  output        io_connPE_41_ready,
  input         io_connPE_41_valid,
  input  [63:0] io_connPE_41_bits,
  output        io_connPE_42_ready,
  input         io_connPE_42_valid,
  input  [63:0] io_connPE_42_bits,
  output        io_connPE_43_ready,
  input         io_connPE_43_valid,
  input  [63:0] io_connPE_43_bits,
  output        io_connPE_44_ready,
  input         io_connPE_44_valid,
  input  [63:0] io_connPE_44_bits,
  output        io_connPE_45_ready,
  input         io_connPE_45_valid,
  input  [63:0] io_connPE_45_bits,
  output        io_connPE_46_ready,
  input         io_connPE_46_valid,
  input  [63:0] io_connPE_46_bits,
  output        io_connPE_47_ready,
  input         io_connPE_47_valid,
  input  [63:0] io_connPE_47_bits,
  output        io_connPE_48_ready,
  input         io_connPE_48_valid,
  input  [63:0] io_connPE_48_bits,
  output        io_connPE_49_ready,
  input         io_connPE_49_valid,
  input  [63:0] io_connPE_49_bits,
  output        io_connPE_50_ready,
  input         io_connPE_50_valid,
  input  [63:0] io_connPE_50_bits,
  output        io_connPE_51_ready,
  input         io_connPE_51_valid,
  input  [63:0] io_connPE_51_bits,
  output        io_connPE_52_ready,
  input         io_connPE_52_valid,
  input  [63:0] io_connPE_52_bits,
  output        io_connPE_53_ready,
  input         io_connPE_53_valid,
  input  [63:0] io_connPE_53_bits,
  output        io_connPE_54_ready,
  input         io_connPE_54_valid,
  input  [63:0] io_connPE_54_bits,
  output        io_connPE_55_ready,
  input         io_connPE_55_valid,
  input  [63:0] io_connPE_55_bits,
  output        io_connPE_56_ready,
  input         io_connPE_56_valid,
  input  [63:0] io_connPE_56_bits,
  output        io_connPE_57_ready,
  input         io_connPE_57_valid,
  input  [63:0] io_connPE_57_bits,
  output        io_connPE_58_ready,
  input         io_connPE_58_valid,
  input  [63:0] io_connPE_58_bits,
  output        io_connPE_59_ready,
  input         io_connPE_59_valid,
  input  [63:0] io_connPE_59_bits,
  output        io_connPE_60_ready,
  input         io_connPE_60_valid,
  input  [63:0] io_connPE_60_bits,
  output        io_connPE_61_ready,
  input         io_connPE_61_valid,
  input  [63:0] io_connPE_61_bits,
  output        io_connPE_62_ready,
  input         io_connPE_62_valid,
  input  [63:0] io_connPE_62_bits,
  output        io_connPE_63_ready,
  input         io_connPE_63_valid,
  input  [63:0] io_connPE_63_bits
);
  wire  networkUnits_0_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_0_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_0_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_0_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_0_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_0_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_0_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_0_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_0_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_0_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_0_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_1_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_1_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_1_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_1_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_1_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_1_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_1_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_1_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_1_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_1_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_1_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_2_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_2_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_2_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_2_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_2_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_2_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_2_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_2_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_2_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_2_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_2_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_3_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_3_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_3_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_3_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_3_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_3_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_3_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_3_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_3_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_3_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_3_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_4_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_4_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_4_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_4_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_4_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_4_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_4_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_4_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_4_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_4_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_4_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_5_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_5_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_5_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_5_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_5_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_5_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_5_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_5_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_5_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_5_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_5_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_6_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_6_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_6_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_6_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_6_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_6_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_6_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_6_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_6_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_6_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_6_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_7_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_7_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_7_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_7_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_7_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_7_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_7_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_7_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_7_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_7_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_7_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_8_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_8_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_8_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_8_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_8_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_8_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_8_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_8_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_8_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_8_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_8_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_9_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_9_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_9_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_9_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_9_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_9_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_9_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_9_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_9_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_9_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_9_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_10_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_10_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_10_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_10_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_10_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_10_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_10_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_10_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_10_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_10_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_10_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_11_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_11_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_11_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_11_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_11_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_11_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_11_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_11_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_11_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_11_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_11_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_12_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_12_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_12_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_12_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_12_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_12_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_12_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_12_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_12_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_12_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_12_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_13_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_13_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_13_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_13_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_13_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_13_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_13_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_13_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_13_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_13_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_13_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_14_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_14_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_14_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_14_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_14_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_14_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_14_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_14_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_14_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_14_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_14_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_15_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_15_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_15_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_15_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_15_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_15_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_15_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_15_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_15_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_15_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_15_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_16_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_16_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_16_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_16_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_16_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_16_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_16_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_16_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_16_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_16_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_16_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_17_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_17_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_17_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_17_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_17_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_17_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_17_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_17_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_17_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_17_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_17_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_18_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_18_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_18_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_18_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_18_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_18_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_18_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_18_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_18_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_18_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_18_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_19_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_19_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_19_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_19_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_19_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_19_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_19_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_19_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_19_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_19_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_19_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_20_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_20_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_20_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_20_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_20_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_20_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_20_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_20_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_20_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_20_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_20_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_21_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_21_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_21_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_21_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_21_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_21_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_21_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_21_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_21_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_21_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_21_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_22_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_22_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_22_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_22_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_22_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_22_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_22_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_22_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_22_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_22_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_22_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_23_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_23_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_23_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_23_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_23_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_23_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_23_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_23_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_23_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_23_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_23_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_24_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_24_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_24_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_24_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_24_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_24_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_24_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_24_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_24_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_24_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_24_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_25_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_25_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_25_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_25_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_25_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_25_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_25_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_25_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_25_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_25_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_25_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_26_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_26_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_26_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_26_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_26_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_26_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_26_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_26_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_26_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_26_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_26_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_27_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_27_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_27_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_27_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_27_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_27_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_27_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_27_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_27_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_27_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_27_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_28_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_28_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_28_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_28_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_28_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_28_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_28_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_28_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_28_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_28_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_28_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_29_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_29_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_29_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_29_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_29_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_29_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_29_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_29_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_29_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_29_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_29_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_30_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_30_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_30_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_30_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_30_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_30_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_30_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_30_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_30_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_30_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_30_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_31_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_31_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_31_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_31_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_31_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_31_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_31_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_31_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_31_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_31_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_31_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_32_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_32_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_32_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_32_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_32_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_32_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_32_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_32_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_32_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_32_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_32_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_33_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_33_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_33_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_33_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_33_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_33_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_33_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_33_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_33_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_33_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_33_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_34_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_34_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_34_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_34_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_34_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_34_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_34_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_34_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_34_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_34_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_34_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_35_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_35_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_35_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_35_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_35_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_35_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_35_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_35_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_35_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_35_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_35_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_36_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_36_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_36_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_36_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_36_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_36_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_36_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_36_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_36_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_36_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_36_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_37_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_37_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_37_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_37_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_37_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_37_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_37_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_37_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_37_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_37_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_37_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_38_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_38_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_38_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_38_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_38_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_38_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_38_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_38_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_38_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_38_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_38_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_39_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_39_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_39_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_39_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_39_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_39_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_39_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_39_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_39_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_39_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_39_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_40_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_40_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_40_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_40_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_40_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_40_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_40_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_40_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_40_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_40_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_40_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_41_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_41_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_41_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_41_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_41_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_41_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_41_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_41_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_41_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_41_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_41_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_42_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_42_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_42_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_42_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_42_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_42_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_42_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_42_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_42_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_42_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_42_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_43_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_43_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_43_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_43_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_43_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_43_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_43_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_43_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_43_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_43_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_43_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_44_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_44_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_44_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_44_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_44_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_44_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_44_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_44_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_44_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_44_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_44_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_45_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_45_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_45_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_45_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_45_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_45_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_45_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_45_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_45_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_45_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_45_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_46_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_46_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_46_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_46_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_46_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_46_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_46_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_46_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_46_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_46_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_46_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_47_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_47_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_47_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_47_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_47_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_47_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_47_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_47_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_47_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_47_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_47_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_48_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_48_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_48_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_48_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_48_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_48_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_48_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_48_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_48_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_48_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_48_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_49_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_49_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_49_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_49_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_49_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_49_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_49_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_49_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_49_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_49_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_49_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_50_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_50_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_50_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_50_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_50_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_50_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_50_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_50_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_50_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_50_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_50_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_51_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_51_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_51_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_51_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_51_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_51_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_51_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_51_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_51_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_51_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_51_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_52_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_52_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_52_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_52_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_52_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_52_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_52_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_52_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_52_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_52_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_52_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_53_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_53_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_53_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_53_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_53_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_53_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_53_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_53_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_53_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_53_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_53_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_54_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_54_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_54_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_54_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_54_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_54_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_54_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_54_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_54_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_54_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_54_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_55_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_55_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_55_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_55_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_55_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_55_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_55_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_55_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_55_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_55_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_55_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_56_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_56_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_56_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_56_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_56_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_56_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_56_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_56_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_56_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_56_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_56_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_57_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_57_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_57_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_57_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_57_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_57_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_57_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_57_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_57_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_57_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_57_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_58_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_58_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_58_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_58_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_58_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_58_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_58_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_58_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_58_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_58_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_58_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_59_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_59_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_59_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_59_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_59_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_59_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_59_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_59_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_59_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_59_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_59_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_60_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_60_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_60_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_60_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_60_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_60_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_60_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_60_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_60_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_60_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_60_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_61_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_61_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_61_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_61_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_61_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_61_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_61_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_61_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_61_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_61_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_61_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_62_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_62_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_62_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_62_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_62_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_62_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_62_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_62_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_62_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_62_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_62_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_63_clock; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_63_reset; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_63_io_addressIn_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_63_io_addressIn_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_63_io_addressIn_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_63_io_peAddress_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_63_io_peAddress_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_63_io_peAddress_bits; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_63_io_addressOut_ready; // @[argRouteNetwork.scala 52:52]
  wire  networkUnits_63_io_addressOut_valid; // @[argRouteNetwork.scala 52:52]
  wire [63:0] networkUnits_63_io_addressOut_bits; // @[argRouteNetwork.scala 52:52]
  wire  virtNetworkUnits_0_clock; // @[argRouteNetwork.scala 67:58]
  wire  virtNetworkUnits_0_reset; // @[argRouteNetwork.scala 67:58]
  wire  virtNetworkUnits_0_io_addressIn_ready; // @[argRouteNetwork.scala 67:58]
  wire  virtNetworkUnits_0_io_addressIn_valid; // @[argRouteNetwork.scala 67:58]
  wire [63:0] virtNetworkUnits_0_io_addressIn_bits; // @[argRouteNetwork.scala 67:58]
  wire  virtNetworkUnits_0_io_vasAddressOut_ready; // @[argRouteNetwork.scala 67:58]
  wire  virtNetworkUnits_0_io_vasAddressOut_valid; // @[argRouteNetwork.scala 67:58]
  wire [63:0] virtNetworkUnits_0_io_vasAddressOut_bits; // @[argRouteNetwork.scala 67:58]
  wire  virtNetworkUnits_1_clock; // @[argRouteNetwork.scala 67:58]
  wire  virtNetworkUnits_1_reset; // @[argRouteNetwork.scala 67:58]
  wire  virtNetworkUnits_1_io_addressIn_ready; // @[argRouteNetwork.scala 67:58]
  wire  virtNetworkUnits_1_io_addressIn_valid; // @[argRouteNetwork.scala 67:58]
  wire [63:0] virtNetworkUnits_1_io_addressIn_bits; // @[argRouteNetwork.scala 67:58]
  wire  virtNetworkUnits_1_io_vasAddressOut_ready; // @[argRouteNetwork.scala 67:58]
  wire  virtNetworkUnits_1_io_vasAddressOut_valid; // @[argRouteNetwork.scala 67:58]
  wire [63:0] virtNetworkUnits_1_io_vasAddressOut_bits; // @[argRouteNetwork.scala 67:58]
  wire  virtNetworkUnits_1_io_addressOut_ready; // @[argRouteNetwork.scala 67:58]
  wire  virtNetworkUnits_1_io_addressOut_valid; // @[argRouteNetwork.scala 67:58]
  wire [63:0] virtNetworkUnits_1_io_addressOut_bits; // @[argRouteNetwork.scala 67:58]
  wire  queues_0_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_0_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_0_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_0_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_0_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_0_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_0_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_0_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_1_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_1_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_1_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_1_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_1_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_1_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_1_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_1_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_2_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_2_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_2_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_2_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_2_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_2_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_2_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_2_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_3_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_3_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_3_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_3_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_3_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_3_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_3_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_3_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_4_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_4_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_4_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_4_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_4_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_4_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_4_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_4_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_5_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_5_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_5_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_5_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_5_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_5_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_5_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_5_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_6_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_6_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_6_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_6_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_6_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_6_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_6_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_6_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_7_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_7_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_7_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_7_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_7_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_7_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_7_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_7_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_8_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_8_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_8_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_8_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_8_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_8_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_8_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_8_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_9_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_9_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_9_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_9_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_9_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_9_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_9_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_9_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_10_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_10_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_10_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_10_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_10_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_10_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_10_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_10_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_11_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_11_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_11_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_11_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_11_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_11_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_11_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_11_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_12_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_12_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_12_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_12_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_12_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_12_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_12_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_12_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_13_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_13_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_13_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_13_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_13_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_13_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_13_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_13_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_14_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_14_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_14_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_14_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_14_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_14_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_14_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_14_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_15_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_15_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_15_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_15_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_15_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_15_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_15_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_15_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_16_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_16_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_16_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_16_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_16_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_16_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_16_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_16_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_17_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_17_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_17_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_17_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_17_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_17_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_17_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_17_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_18_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_18_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_18_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_18_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_18_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_18_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_18_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_18_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_19_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_19_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_19_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_19_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_19_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_19_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_19_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_19_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_20_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_20_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_20_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_20_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_20_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_20_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_20_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_20_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_21_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_21_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_21_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_21_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_21_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_21_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_21_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_21_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_22_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_22_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_22_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_22_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_22_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_22_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_22_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_22_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_23_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_23_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_23_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_23_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_23_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_23_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_23_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_23_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_24_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_24_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_24_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_24_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_24_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_24_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_24_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_24_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_25_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_25_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_25_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_25_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_25_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_25_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_25_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_25_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_26_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_26_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_26_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_26_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_26_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_26_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_26_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_26_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_27_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_27_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_27_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_27_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_27_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_27_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_27_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_27_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_28_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_28_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_28_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_28_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_28_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_28_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_28_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_28_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_29_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_29_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_29_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_29_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_29_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_29_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_29_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_29_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_30_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_30_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_30_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_30_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_30_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_30_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_30_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_30_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_31_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_31_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_31_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_31_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_31_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_31_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_31_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_31_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_32_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_32_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_32_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_32_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_32_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_32_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_32_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_32_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_33_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_33_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_33_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_33_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_33_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_33_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_33_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_33_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_34_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_34_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_34_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_34_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_34_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_34_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_34_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_34_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_35_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_35_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_35_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_35_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_35_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_35_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_35_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_35_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_36_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_36_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_36_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_36_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_36_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_36_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_36_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_36_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_37_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_37_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_37_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_37_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_37_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_37_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_37_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_37_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_38_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_38_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_38_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_38_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_38_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_38_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_38_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_38_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_39_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_39_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_39_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_39_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_39_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_39_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_39_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_39_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_40_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_40_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_40_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_40_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_40_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_40_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_40_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_40_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_41_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_41_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_41_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_41_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_41_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_41_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_41_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_41_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_42_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_42_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_42_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_42_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_42_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_42_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_42_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_42_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_43_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_43_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_43_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_43_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_43_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_43_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_43_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_43_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_44_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_44_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_44_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_44_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_44_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_44_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_44_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_44_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_45_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_45_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_45_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_45_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_45_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_45_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_45_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_45_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_46_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_46_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_46_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_46_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_46_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_46_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_46_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_46_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_47_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_47_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_47_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_47_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_47_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_47_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_47_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_47_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_48_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_48_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_48_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_48_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_48_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_48_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_48_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_48_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_49_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_49_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_49_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_49_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_49_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_49_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_49_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_49_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_50_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_50_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_50_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_50_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_50_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_50_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_50_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_50_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_51_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_51_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_51_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_51_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_51_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_51_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_51_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_51_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_52_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_52_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_52_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_52_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_52_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_52_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_52_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_52_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_53_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_53_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_53_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_53_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_53_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_53_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_53_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_53_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_54_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_54_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_54_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_54_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_54_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_54_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_54_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_54_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_55_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_55_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_55_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_55_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_55_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_55_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_55_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_55_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_56_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_56_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_56_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_56_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_56_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_56_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_56_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_56_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_57_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_57_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_57_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_57_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_57_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_57_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_57_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_57_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_58_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_58_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_58_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_58_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_58_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_58_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_58_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_58_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_59_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_59_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_59_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_59_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_59_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_59_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_59_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_59_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_60_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_60_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_60_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_60_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_60_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_60_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_60_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_60_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_61_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_61_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_61_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_61_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_61_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_61_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_61_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_61_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_62_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_62_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_62_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_62_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_62_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_62_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_62_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_62_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_63_clock; // @[argRouteNetwork.scala 79:49]
  wire  queues_63_reset; // @[argRouteNetwork.scala 79:49]
  wire  queues_63_io_addressIn_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_63_io_addressIn_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_63_io_addressIn_bits; // @[argRouteNetwork.scala 79:49]
  wire  queues_63_io_addressOut_ready; // @[argRouteNetwork.scala 79:49]
  wire  queues_63_io_addressOut_valid; // @[argRouteNetwork.scala 79:49]
  wire [63:0] queues_63_io_addressOut_bits; // @[argRouteNetwork.scala 79:49]
  argRouteNtwUnit networkUnits_0 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_0_clock),
    .reset(networkUnits_0_reset),
    .io_addressIn_ready(networkUnits_0_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_0_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_0_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_0_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_0_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_0_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_0_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_0_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_0_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_1 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_1_clock),
    .reset(networkUnits_1_reset),
    .io_addressIn_ready(networkUnits_1_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_1_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_1_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_1_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_1_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_1_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_1_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_1_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_1_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_2 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_2_clock),
    .reset(networkUnits_2_reset),
    .io_addressIn_ready(networkUnits_2_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_2_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_2_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_2_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_2_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_2_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_2_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_2_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_2_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_3 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_3_clock),
    .reset(networkUnits_3_reset),
    .io_addressIn_ready(networkUnits_3_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_3_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_3_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_3_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_3_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_3_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_3_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_3_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_3_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_4 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_4_clock),
    .reset(networkUnits_4_reset),
    .io_addressIn_ready(networkUnits_4_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_4_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_4_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_4_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_4_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_4_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_4_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_4_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_4_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_5 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_5_clock),
    .reset(networkUnits_5_reset),
    .io_addressIn_ready(networkUnits_5_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_5_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_5_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_5_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_5_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_5_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_5_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_5_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_5_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_6 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_6_clock),
    .reset(networkUnits_6_reset),
    .io_addressIn_ready(networkUnits_6_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_6_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_6_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_6_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_6_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_6_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_6_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_6_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_6_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_7 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_7_clock),
    .reset(networkUnits_7_reset),
    .io_addressIn_ready(networkUnits_7_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_7_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_7_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_7_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_7_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_7_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_7_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_7_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_7_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_8 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_8_clock),
    .reset(networkUnits_8_reset),
    .io_addressIn_ready(networkUnits_8_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_8_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_8_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_8_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_8_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_8_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_8_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_8_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_8_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_9 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_9_clock),
    .reset(networkUnits_9_reset),
    .io_addressIn_ready(networkUnits_9_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_9_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_9_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_9_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_9_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_9_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_9_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_9_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_9_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_10 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_10_clock),
    .reset(networkUnits_10_reset),
    .io_addressIn_ready(networkUnits_10_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_10_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_10_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_10_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_10_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_10_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_10_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_10_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_10_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_11 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_11_clock),
    .reset(networkUnits_11_reset),
    .io_addressIn_ready(networkUnits_11_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_11_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_11_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_11_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_11_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_11_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_11_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_11_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_11_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_12 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_12_clock),
    .reset(networkUnits_12_reset),
    .io_addressIn_ready(networkUnits_12_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_12_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_12_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_12_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_12_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_12_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_12_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_12_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_12_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_13 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_13_clock),
    .reset(networkUnits_13_reset),
    .io_addressIn_ready(networkUnits_13_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_13_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_13_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_13_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_13_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_13_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_13_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_13_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_13_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_14 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_14_clock),
    .reset(networkUnits_14_reset),
    .io_addressIn_ready(networkUnits_14_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_14_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_14_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_14_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_14_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_14_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_14_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_14_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_14_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_15 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_15_clock),
    .reset(networkUnits_15_reset),
    .io_addressIn_ready(networkUnits_15_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_15_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_15_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_15_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_15_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_15_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_15_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_15_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_15_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_16 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_16_clock),
    .reset(networkUnits_16_reset),
    .io_addressIn_ready(networkUnits_16_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_16_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_16_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_16_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_16_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_16_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_16_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_16_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_16_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_17 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_17_clock),
    .reset(networkUnits_17_reset),
    .io_addressIn_ready(networkUnits_17_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_17_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_17_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_17_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_17_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_17_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_17_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_17_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_17_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_18 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_18_clock),
    .reset(networkUnits_18_reset),
    .io_addressIn_ready(networkUnits_18_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_18_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_18_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_18_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_18_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_18_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_18_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_18_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_18_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_19 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_19_clock),
    .reset(networkUnits_19_reset),
    .io_addressIn_ready(networkUnits_19_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_19_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_19_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_19_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_19_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_19_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_19_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_19_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_19_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_20 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_20_clock),
    .reset(networkUnits_20_reset),
    .io_addressIn_ready(networkUnits_20_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_20_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_20_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_20_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_20_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_20_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_20_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_20_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_20_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_21 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_21_clock),
    .reset(networkUnits_21_reset),
    .io_addressIn_ready(networkUnits_21_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_21_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_21_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_21_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_21_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_21_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_21_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_21_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_21_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_22 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_22_clock),
    .reset(networkUnits_22_reset),
    .io_addressIn_ready(networkUnits_22_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_22_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_22_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_22_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_22_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_22_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_22_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_22_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_22_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_23 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_23_clock),
    .reset(networkUnits_23_reset),
    .io_addressIn_ready(networkUnits_23_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_23_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_23_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_23_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_23_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_23_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_23_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_23_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_23_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_24 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_24_clock),
    .reset(networkUnits_24_reset),
    .io_addressIn_ready(networkUnits_24_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_24_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_24_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_24_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_24_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_24_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_24_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_24_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_24_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_25 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_25_clock),
    .reset(networkUnits_25_reset),
    .io_addressIn_ready(networkUnits_25_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_25_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_25_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_25_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_25_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_25_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_25_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_25_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_25_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_26 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_26_clock),
    .reset(networkUnits_26_reset),
    .io_addressIn_ready(networkUnits_26_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_26_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_26_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_26_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_26_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_26_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_26_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_26_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_26_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_27 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_27_clock),
    .reset(networkUnits_27_reset),
    .io_addressIn_ready(networkUnits_27_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_27_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_27_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_27_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_27_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_27_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_27_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_27_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_27_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_28 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_28_clock),
    .reset(networkUnits_28_reset),
    .io_addressIn_ready(networkUnits_28_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_28_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_28_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_28_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_28_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_28_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_28_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_28_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_28_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_29 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_29_clock),
    .reset(networkUnits_29_reset),
    .io_addressIn_ready(networkUnits_29_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_29_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_29_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_29_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_29_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_29_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_29_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_29_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_29_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_30 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_30_clock),
    .reset(networkUnits_30_reset),
    .io_addressIn_ready(networkUnits_30_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_30_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_30_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_30_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_30_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_30_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_30_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_30_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_30_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_31 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_31_clock),
    .reset(networkUnits_31_reset),
    .io_addressIn_ready(networkUnits_31_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_31_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_31_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_31_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_31_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_31_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_31_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_31_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_31_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_32 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_32_clock),
    .reset(networkUnits_32_reset),
    .io_addressIn_ready(networkUnits_32_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_32_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_32_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_32_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_32_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_32_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_32_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_32_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_32_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_33 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_33_clock),
    .reset(networkUnits_33_reset),
    .io_addressIn_ready(networkUnits_33_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_33_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_33_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_33_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_33_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_33_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_33_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_33_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_33_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_34 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_34_clock),
    .reset(networkUnits_34_reset),
    .io_addressIn_ready(networkUnits_34_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_34_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_34_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_34_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_34_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_34_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_34_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_34_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_34_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_35 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_35_clock),
    .reset(networkUnits_35_reset),
    .io_addressIn_ready(networkUnits_35_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_35_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_35_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_35_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_35_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_35_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_35_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_35_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_35_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_36 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_36_clock),
    .reset(networkUnits_36_reset),
    .io_addressIn_ready(networkUnits_36_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_36_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_36_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_36_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_36_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_36_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_36_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_36_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_36_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_37 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_37_clock),
    .reset(networkUnits_37_reset),
    .io_addressIn_ready(networkUnits_37_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_37_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_37_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_37_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_37_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_37_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_37_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_37_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_37_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_38 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_38_clock),
    .reset(networkUnits_38_reset),
    .io_addressIn_ready(networkUnits_38_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_38_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_38_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_38_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_38_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_38_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_38_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_38_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_38_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_39 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_39_clock),
    .reset(networkUnits_39_reset),
    .io_addressIn_ready(networkUnits_39_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_39_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_39_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_39_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_39_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_39_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_39_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_39_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_39_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_40 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_40_clock),
    .reset(networkUnits_40_reset),
    .io_addressIn_ready(networkUnits_40_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_40_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_40_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_40_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_40_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_40_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_40_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_40_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_40_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_41 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_41_clock),
    .reset(networkUnits_41_reset),
    .io_addressIn_ready(networkUnits_41_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_41_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_41_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_41_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_41_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_41_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_41_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_41_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_41_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_42 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_42_clock),
    .reset(networkUnits_42_reset),
    .io_addressIn_ready(networkUnits_42_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_42_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_42_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_42_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_42_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_42_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_42_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_42_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_42_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_43 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_43_clock),
    .reset(networkUnits_43_reset),
    .io_addressIn_ready(networkUnits_43_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_43_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_43_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_43_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_43_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_43_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_43_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_43_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_43_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_44 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_44_clock),
    .reset(networkUnits_44_reset),
    .io_addressIn_ready(networkUnits_44_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_44_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_44_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_44_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_44_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_44_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_44_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_44_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_44_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_45 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_45_clock),
    .reset(networkUnits_45_reset),
    .io_addressIn_ready(networkUnits_45_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_45_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_45_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_45_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_45_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_45_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_45_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_45_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_45_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_46 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_46_clock),
    .reset(networkUnits_46_reset),
    .io_addressIn_ready(networkUnits_46_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_46_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_46_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_46_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_46_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_46_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_46_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_46_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_46_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_47 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_47_clock),
    .reset(networkUnits_47_reset),
    .io_addressIn_ready(networkUnits_47_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_47_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_47_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_47_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_47_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_47_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_47_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_47_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_47_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_48 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_48_clock),
    .reset(networkUnits_48_reset),
    .io_addressIn_ready(networkUnits_48_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_48_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_48_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_48_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_48_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_48_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_48_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_48_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_48_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_49 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_49_clock),
    .reset(networkUnits_49_reset),
    .io_addressIn_ready(networkUnits_49_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_49_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_49_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_49_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_49_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_49_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_49_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_49_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_49_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_50 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_50_clock),
    .reset(networkUnits_50_reset),
    .io_addressIn_ready(networkUnits_50_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_50_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_50_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_50_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_50_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_50_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_50_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_50_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_50_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_51 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_51_clock),
    .reset(networkUnits_51_reset),
    .io_addressIn_ready(networkUnits_51_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_51_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_51_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_51_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_51_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_51_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_51_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_51_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_51_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_52 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_52_clock),
    .reset(networkUnits_52_reset),
    .io_addressIn_ready(networkUnits_52_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_52_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_52_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_52_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_52_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_52_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_52_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_52_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_52_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_53 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_53_clock),
    .reset(networkUnits_53_reset),
    .io_addressIn_ready(networkUnits_53_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_53_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_53_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_53_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_53_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_53_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_53_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_53_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_53_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_54 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_54_clock),
    .reset(networkUnits_54_reset),
    .io_addressIn_ready(networkUnits_54_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_54_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_54_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_54_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_54_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_54_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_54_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_54_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_54_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_55 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_55_clock),
    .reset(networkUnits_55_reset),
    .io_addressIn_ready(networkUnits_55_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_55_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_55_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_55_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_55_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_55_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_55_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_55_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_55_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_56 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_56_clock),
    .reset(networkUnits_56_reset),
    .io_addressIn_ready(networkUnits_56_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_56_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_56_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_56_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_56_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_56_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_56_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_56_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_56_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_57 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_57_clock),
    .reset(networkUnits_57_reset),
    .io_addressIn_ready(networkUnits_57_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_57_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_57_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_57_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_57_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_57_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_57_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_57_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_57_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_58 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_58_clock),
    .reset(networkUnits_58_reset),
    .io_addressIn_ready(networkUnits_58_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_58_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_58_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_58_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_58_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_58_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_58_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_58_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_58_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_59 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_59_clock),
    .reset(networkUnits_59_reset),
    .io_addressIn_ready(networkUnits_59_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_59_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_59_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_59_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_59_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_59_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_59_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_59_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_59_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_60 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_60_clock),
    .reset(networkUnits_60_reset),
    .io_addressIn_ready(networkUnits_60_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_60_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_60_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_60_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_60_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_60_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_60_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_60_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_60_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_61 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_61_clock),
    .reset(networkUnits_61_reset),
    .io_addressIn_ready(networkUnits_61_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_61_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_61_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_61_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_61_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_61_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_61_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_61_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_61_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_62 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_62_clock),
    .reset(networkUnits_62_reset),
    .io_addressIn_ready(networkUnits_62_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_62_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_62_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_62_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_62_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_62_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_62_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_62_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_62_io_addressOut_bits)
  );
  argRouteNtwUnit networkUnits_63 ( // @[argRouteNetwork.scala 52:52]
    .clock(networkUnits_63_clock),
    .reset(networkUnits_63_reset),
    .io_addressIn_ready(networkUnits_63_io_addressIn_ready),
    .io_addressIn_valid(networkUnits_63_io_addressIn_valid),
    .io_addressIn_bits(networkUnits_63_io_addressIn_bits),
    .io_peAddress_ready(networkUnits_63_io_peAddress_ready),
    .io_peAddress_valid(networkUnits_63_io_peAddress_valid),
    .io_peAddress_bits(networkUnits_63_io_peAddress_bits),
    .io_addressOut_ready(networkUnits_63_io_addressOut_ready),
    .io_addressOut_valid(networkUnits_63_io_addressOut_valid),
    .io_addressOut_bits(networkUnits_63_io_addressOut_bits)
  );
  argRouteNtwVirtUnit virtNetworkUnits_0 ( // @[argRouteNetwork.scala 67:58]
    .clock(virtNetworkUnits_0_clock),
    .reset(virtNetworkUnits_0_reset),
    .io_addressIn_ready(virtNetworkUnits_0_io_addressIn_ready),
    .io_addressIn_valid(virtNetworkUnits_0_io_addressIn_valid),
    .io_addressIn_bits(virtNetworkUnits_0_io_addressIn_bits),
    .io_vasAddressOut_ready(virtNetworkUnits_0_io_vasAddressOut_ready),
    .io_vasAddressOut_valid(virtNetworkUnits_0_io_vasAddressOut_valid),
    .io_vasAddressOut_bits(virtNetworkUnits_0_io_vasAddressOut_bits)
  );
  argRouteNtwVirtUnit_1 virtNetworkUnits_1 ( // @[argRouteNetwork.scala 67:58]
    .clock(virtNetworkUnits_1_clock),
    .reset(virtNetworkUnits_1_reset),
    .io_addressIn_ready(virtNetworkUnits_1_io_addressIn_ready),
    .io_addressIn_valid(virtNetworkUnits_1_io_addressIn_valid),
    .io_addressIn_bits(virtNetworkUnits_1_io_addressIn_bits),
    .io_vasAddressOut_ready(virtNetworkUnits_1_io_vasAddressOut_ready),
    .io_vasAddressOut_valid(virtNetworkUnits_1_io_vasAddressOut_valid),
    .io_vasAddressOut_bits(virtNetworkUnits_1_io_vasAddressOut_bits),
    .io_addressOut_ready(virtNetworkUnits_1_io_addressOut_ready),
    .io_addressOut_valid(virtNetworkUnits_1_io_addressOut_valid),
    .io_addressOut_bits(virtNetworkUnits_1_io_addressOut_bits)
  );
  contQueue_64 queues_0 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_0_clock),
    .reset(queues_0_reset),
    .io_addressIn_ready(queues_0_io_addressIn_ready),
    .io_addressIn_valid(queues_0_io_addressIn_valid),
    .io_addressIn_bits(queues_0_io_addressIn_bits),
    .io_addressOut_ready(queues_0_io_addressOut_ready),
    .io_addressOut_valid(queues_0_io_addressOut_valid),
    .io_addressOut_bits(queues_0_io_addressOut_bits)
  );
  contQueue_64 queues_1 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_1_clock),
    .reset(queues_1_reset),
    .io_addressIn_ready(queues_1_io_addressIn_ready),
    .io_addressIn_valid(queues_1_io_addressIn_valid),
    .io_addressIn_bits(queues_1_io_addressIn_bits),
    .io_addressOut_ready(queues_1_io_addressOut_ready),
    .io_addressOut_valid(queues_1_io_addressOut_valid),
    .io_addressOut_bits(queues_1_io_addressOut_bits)
  );
  contQueue_64 queues_2 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_2_clock),
    .reset(queues_2_reset),
    .io_addressIn_ready(queues_2_io_addressIn_ready),
    .io_addressIn_valid(queues_2_io_addressIn_valid),
    .io_addressIn_bits(queues_2_io_addressIn_bits),
    .io_addressOut_ready(queues_2_io_addressOut_ready),
    .io_addressOut_valid(queues_2_io_addressOut_valid),
    .io_addressOut_bits(queues_2_io_addressOut_bits)
  );
  contQueue_64 queues_3 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_3_clock),
    .reset(queues_3_reset),
    .io_addressIn_ready(queues_3_io_addressIn_ready),
    .io_addressIn_valid(queues_3_io_addressIn_valid),
    .io_addressIn_bits(queues_3_io_addressIn_bits),
    .io_addressOut_ready(queues_3_io_addressOut_ready),
    .io_addressOut_valid(queues_3_io_addressOut_valid),
    .io_addressOut_bits(queues_3_io_addressOut_bits)
  );
  contQueue_64 queues_4 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_4_clock),
    .reset(queues_4_reset),
    .io_addressIn_ready(queues_4_io_addressIn_ready),
    .io_addressIn_valid(queues_4_io_addressIn_valid),
    .io_addressIn_bits(queues_4_io_addressIn_bits),
    .io_addressOut_ready(queues_4_io_addressOut_ready),
    .io_addressOut_valid(queues_4_io_addressOut_valid),
    .io_addressOut_bits(queues_4_io_addressOut_bits)
  );
  contQueue_64 queues_5 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_5_clock),
    .reset(queues_5_reset),
    .io_addressIn_ready(queues_5_io_addressIn_ready),
    .io_addressIn_valid(queues_5_io_addressIn_valid),
    .io_addressIn_bits(queues_5_io_addressIn_bits),
    .io_addressOut_ready(queues_5_io_addressOut_ready),
    .io_addressOut_valid(queues_5_io_addressOut_valid),
    .io_addressOut_bits(queues_5_io_addressOut_bits)
  );
  contQueue_64 queues_6 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_6_clock),
    .reset(queues_6_reset),
    .io_addressIn_ready(queues_6_io_addressIn_ready),
    .io_addressIn_valid(queues_6_io_addressIn_valid),
    .io_addressIn_bits(queues_6_io_addressIn_bits),
    .io_addressOut_ready(queues_6_io_addressOut_ready),
    .io_addressOut_valid(queues_6_io_addressOut_valid),
    .io_addressOut_bits(queues_6_io_addressOut_bits)
  );
  contQueue_64 queues_7 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_7_clock),
    .reset(queues_7_reset),
    .io_addressIn_ready(queues_7_io_addressIn_ready),
    .io_addressIn_valid(queues_7_io_addressIn_valid),
    .io_addressIn_bits(queues_7_io_addressIn_bits),
    .io_addressOut_ready(queues_7_io_addressOut_ready),
    .io_addressOut_valid(queues_7_io_addressOut_valid),
    .io_addressOut_bits(queues_7_io_addressOut_bits)
  );
  contQueue_64 queues_8 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_8_clock),
    .reset(queues_8_reset),
    .io_addressIn_ready(queues_8_io_addressIn_ready),
    .io_addressIn_valid(queues_8_io_addressIn_valid),
    .io_addressIn_bits(queues_8_io_addressIn_bits),
    .io_addressOut_ready(queues_8_io_addressOut_ready),
    .io_addressOut_valid(queues_8_io_addressOut_valid),
    .io_addressOut_bits(queues_8_io_addressOut_bits)
  );
  contQueue_64 queues_9 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_9_clock),
    .reset(queues_9_reset),
    .io_addressIn_ready(queues_9_io_addressIn_ready),
    .io_addressIn_valid(queues_9_io_addressIn_valid),
    .io_addressIn_bits(queues_9_io_addressIn_bits),
    .io_addressOut_ready(queues_9_io_addressOut_ready),
    .io_addressOut_valid(queues_9_io_addressOut_valid),
    .io_addressOut_bits(queues_9_io_addressOut_bits)
  );
  contQueue_64 queues_10 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_10_clock),
    .reset(queues_10_reset),
    .io_addressIn_ready(queues_10_io_addressIn_ready),
    .io_addressIn_valid(queues_10_io_addressIn_valid),
    .io_addressIn_bits(queues_10_io_addressIn_bits),
    .io_addressOut_ready(queues_10_io_addressOut_ready),
    .io_addressOut_valid(queues_10_io_addressOut_valid),
    .io_addressOut_bits(queues_10_io_addressOut_bits)
  );
  contQueue_64 queues_11 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_11_clock),
    .reset(queues_11_reset),
    .io_addressIn_ready(queues_11_io_addressIn_ready),
    .io_addressIn_valid(queues_11_io_addressIn_valid),
    .io_addressIn_bits(queues_11_io_addressIn_bits),
    .io_addressOut_ready(queues_11_io_addressOut_ready),
    .io_addressOut_valid(queues_11_io_addressOut_valid),
    .io_addressOut_bits(queues_11_io_addressOut_bits)
  );
  contQueue_64 queues_12 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_12_clock),
    .reset(queues_12_reset),
    .io_addressIn_ready(queues_12_io_addressIn_ready),
    .io_addressIn_valid(queues_12_io_addressIn_valid),
    .io_addressIn_bits(queues_12_io_addressIn_bits),
    .io_addressOut_ready(queues_12_io_addressOut_ready),
    .io_addressOut_valid(queues_12_io_addressOut_valid),
    .io_addressOut_bits(queues_12_io_addressOut_bits)
  );
  contQueue_64 queues_13 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_13_clock),
    .reset(queues_13_reset),
    .io_addressIn_ready(queues_13_io_addressIn_ready),
    .io_addressIn_valid(queues_13_io_addressIn_valid),
    .io_addressIn_bits(queues_13_io_addressIn_bits),
    .io_addressOut_ready(queues_13_io_addressOut_ready),
    .io_addressOut_valid(queues_13_io_addressOut_valid),
    .io_addressOut_bits(queues_13_io_addressOut_bits)
  );
  contQueue_64 queues_14 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_14_clock),
    .reset(queues_14_reset),
    .io_addressIn_ready(queues_14_io_addressIn_ready),
    .io_addressIn_valid(queues_14_io_addressIn_valid),
    .io_addressIn_bits(queues_14_io_addressIn_bits),
    .io_addressOut_ready(queues_14_io_addressOut_ready),
    .io_addressOut_valid(queues_14_io_addressOut_valid),
    .io_addressOut_bits(queues_14_io_addressOut_bits)
  );
  contQueue_64 queues_15 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_15_clock),
    .reset(queues_15_reset),
    .io_addressIn_ready(queues_15_io_addressIn_ready),
    .io_addressIn_valid(queues_15_io_addressIn_valid),
    .io_addressIn_bits(queues_15_io_addressIn_bits),
    .io_addressOut_ready(queues_15_io_addressOut_ready),
    .io_addressOut_valid(queues_15_io_addressOut_valid),
    .io_addressOut_bits(queues_15_io_addressOut_bits)
  );
  contQueue_64 queues_16 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_16_clock),
    .reset(queues_16_reset),
    .io_addressIn_ready(queues_16_io_addressIn_ready),
    .io_addressIn_valid(queues_16_io_addressIn_valid),
    .io_addressIn_bits(queues_16_io_addressIn_bits),
    .io_addressOut_ready(queues_16_io_addressOut_ready),
    .io_addressOut_valid(queues_16_io_addressOut_valid),
    .io_addressOut_bits(queues_16_io_addressOut_bits)
  );
  contQueue_64 queues_17 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_17_clock),
    .reset(queues_17_reset),
    .io_addressIn_ready(queues_17_io_addressIn_ready),
    .io_addressIn_valid(queues_17_io_addressIn_valid),
    .io_addressIn_bits(queues_17_io_addressIn_bits),
    .io_addressOut_ready(queues_17_io_addressOut_ready),
    .io_addressOut_valid(queues_17_io_addressOut_valid),
    .io_addressOut_bits(queues_17_io_addressOut_bits)
  );
  contQueue_64 queues_18 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_18_clock),
    .reset(queues_18_reset),
    .io_addressIn_ready(queues_18_io_addressIn_ready),
    .io_addressIn_valid(queues_18_io_addressIn_valid),
    .io_addressIn_bits(queues_18_io_addressIn_bits),
    .io_addressOut_ready(queues_18_io_addressOut_ready),
    .io_addressOut_valid(queues_18_io_addressOut_valid),
    .io_addressOut_bits(queues_18_io_addressOut_bits)
  );
  contQueue_64 queues_19 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_19_clock),
    .reset(queues_19_reset),
    .io_addressIn_ready(queues_19_io_addressIn_ready),
    .io_addressIn_valid(queues_19_io_addressIn_valid),
    .io_addressIn_bits(queues_19_io_addressIn_bits),
    .io_addressOut_ready(queues_19_io_addressOut_ready),
    .io_addressOut_valid(queues_19_io_addressOut_valid),
    .io_addressOut_bits(queues_19_io_addressOut_bits)
  );
  contQueue_64 queues_20 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_20_clock),
    .reset(queues_20_reset),
    .io_addressIn_ready(queues_20_io_addressIn_ready),
    .io_addressIn_valid(queues_20_io_addressIn_valid),
    .io_addressIn_bits(queues_20_io_addressIn_bits),
    .io_addressOut_ready(queues_20_io_addressOut_ready),
    .io_addressOut_valid(queues_20_io_addressOut_valid),
    .io_addressOut_bits(queues_20_io_addressOut_bits)
  );
  contQueue_64 queues_21 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_21_clock),
    .reset(queues_21_reset),
    .io_addressIn_ready(queues_21_io_addressIn_ready),
    .io_addressIn_valid(queues_21_io_addressIn_valid),
    .io_addressIn_bits(queues_21_io_addressIn_bits),
    .io_addressOut_ready(queues_21_io_addressOut_ready),
    .io_addressOut_valid(queues_21_io_addressOut_valid),
    .io_addressOut_bits(queues_21_io_addressOut_bits)
  );
  contQueue_64 queues_22 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_22_clock),
    .reset(queues_22_reset),
    .io_addressIn_ready(queues_22_io_addressIn_ready),
    .io_addressIn_valid(queues_22_io_addressIn_valid),
    .io_addressIn_bits(queues_22_io_addressIn_bits),
    .io_addressOut_ready(queues_22_io_addressOut_ready),
    .io_addressOut_valid(queues_22_io_addressOut_valid),
    .io_addressOut_bits(queues_22_io_addressOut_bits)
  );
  contQueue_64 queues_23 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_23_clock),
    .reset(queues_23_reset),
    .io_addressIn_ready(queues_23_io_addressIn_ready),
    .io_addressIn_valid(queues_23_io_addressIn_valid),
    .io_addressIn_bits(queues_23_io_addressIn_bits),
    .io_addressOut_ready(queues_23_io_addressOut_ready),
    .io_addressOut_valid(queues_23_io_addressOut_valid),
    .io_addressOut_bits(queues_23_io_addressOut_bits)
  );
  contQueue_64 queues_24 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_24_clock),
    .reset(queues_24_reset),
    .io_addressIn_ready(queues_24_io_addressIn_ready),
    .io_addressIn_valid(queues_24_io_addressIn_valid),
    .io_addressIn_bits(queues_24_io_addressIn_bits),
    .io_addressOut_ready(queues_24_io_addressOut_ready),
    .io_addressOut_valid(queues_24_io_addressOut_valid),
    .io_addressOut_bits(queues_24_io_addressOut_bits)
  );
  contQueue_64 queues_25 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_25_clock),
    .reset(queues_25_reset),
    .io_addressIn_ready(queues_25_io_addressIn_ready),
    .io_addressIn_valid(queues_25_io_addressIn_valid),
    .io_addressIn_bits(queues_25_io_addressIn_bits),
    .io_addressOut_ready(queues_25_io_addressOut_ready),
    .io_addressOut_valid(queues_25_io_addressOut_valid),
    .io_addressOut_bits(queues_25_io_addressOut_bits)
  );
  contQueue_64 queues_26 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_26_clock),
    .reset(queues_26_reset),
    .io_addressIn_ready(queues_26_io_addressIn_ready),
    .io_addressIn_valid(queues_26_io_addressIn_valid),
    .io_addressIn_bits(queues_26_io_addressIn_bits),
    .io_addressOut_ready(queues_26_io_addressOut_ready),
    .io_addressOut_valid(queues_26_io_addressOut_valid),
    .io_addressOut_bits(queues_26_io_addressOut_bits)
  );
  contQueue_64 queues_27 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_27_clock),
    .reset(queues_27_reset),
    .io_addressIn_ready(queues_27_io_addressIn_ready),
    .io_addressIn_valid(queues_27_io_addressIn_valid),
    .io_addressIn_bits(queues_27_io_addressIn_bits),
    .io_addressOut_ready(queues_27_io_addressOut_ready),
    .io_addressOut_valid(queues_27_io_addressOut_valid),
    .io_addressOut_bits(queues_27_io_addressOut_bits)
  );
  contQueue_64 queues_28 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_28_clock),
    .reset(queues_28_reset),
    .io_addressIn_ready(queues_28_io_addressIn_ready),
    .io_addressIn_valid(queues_28_io_addressIn_valid),
    .io_addressIn_bits(queues_28_io_addressIn_bits),
    .io_addressOut_ready(queues_28_io_addressOut_ready),
    .io_addressOut_valid(queues_28_io_addressOut_valid),
    .io_addressOut_bits(queues_28_io_addressOut_bits)
  );
  contQueue_64 queues_29 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_29_clock),
    .reset(queues_29_reset),
    .io_addressIn_ready(queues_29_io_addressIn_ready),
    .io_addressIn_valid(queues_29_io_addressIn_valid),
    .io_addressIn_bits(queues_29_io_addressIn_bits),
    .io_addressOut_ready(queues_29_io_addressOut_ready),
    .io_addressOut_valid(queues_29_io_addressOut_valid),
    .io_addressOut_bits(queues_29_io_addressOut_bits)
  );
  contQueue_64 queues_30 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_30_clock),
    .reset(queues_30_reset),
    .io_addressIn_ready(queues_30_io_addressIn_ready),
    .io_addressIn_valid(queues_30_io_addressIn_valid),
    .io_addressIn_bits(queues_30_io_addressIn_bits),
    .io_addressOut_ready(queues_30_io_addressOut_ready),
    .io_addressOut_valid(queues_30_io_addressOut_valid),
    .io_addressOut_bits(queues_30_io_addressOut_bits)
  );
  contQueue_64 queues_31 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_31_clock),
    .reset(queues_31_reset),
    .io_addressIn_ready(queues_31_io_addressIn_ready),
    .io_addressIn_valid(queues_31_io_addressIn_valid),
    .io_addressIn_bits(queues_31_io_addressIn_bits),
    .io_addressOut_ready(queues_31_io_addressOut_ready),
    .io_addressOut_valid(queues_31_io_addressOut_valid),
    .io_addressOut_bits(queues_31_io_addressOut_bits)
  );
  contQueue_64 queues_32 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_32_clock),
    .reset(queues_32_reset),
    .io_addressIn_ready(queues_32_io_addressIn_ready),
    .io_addressIn_valid(queues_32_io_addressIn_valid),
    .io_addressIn_bits(queues_32_io_addressIn_bits),
    .io_addressOut_ready(queues_32_io_addressOut_ready),
    .io_addressOut_valid(queues_32_io_addressOut_valid),
    .io_addressOut_bits(queues_32_io_addressOut_bits)
  );
  contQueue_64 queues_33 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_33_clock),
    .reset(queues_33_reset),
    .io_addressIn_ready(queues_33_io_addressIn_ready),
    .io_addressIn_valid(queues_33_io_addressIn_valid),
    .io_addressIn_bits(queues_33_io_addressIn_bits),
    .io_addressOut_ready(queues_33_io_addressOut_ready),
    .io_addressOut_valid(queues_33_io_addressOut_valid),
    .io_addressOut_bits(queues_33_io_addressOut_bits)
  );
  contQueue_64 queues_34 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_34_clock),
    .reset(queues_34_reset),
    .io_addressIn_ready(queues_34_io_addressIn_ready),
    .io_addressIn_valid(queues_34_io_addressIn_valid),
    .io_addressIn_bits(queues_34_io_addressIn_bits),
    .io_addressOut_ready(queues_34_io_addressOut_ready),
    .io_addressOut_valid(queues_34_io_addressOut_valid),
    .io_addressOut_bits(queues_34_io_addressOut_bits)
  );
  contQueue_64 queues_35 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_35_clock),
    .reset(queues_35_reset),
    .io_addressIn_ready(queues_35_io_addressIn_ready),
    .io_addressIn_valid(queues_35_io_addressIn_valid),
    .io_addressIn_bits(queues_35_io_addressIn_bits),
    .io_addressOut_ready(queues_35_io_addressOut_ready),
    .io_addressOut_valid(queues_35_io_addressOut_valid),
    .io_addressOut_bits(queues_35_io_addressOut_bits)
  );
  contQueue_64 queues_36 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_36_clock),
    .reset(queues_36_reset),
    .io_addressIn_ready(queues_36_io_addressIn_ready),
    .io_addressIn_valid(queues_36_io_addressIn_valid),
    .io_addressIn_bits(queues_36_io_addressIn_bits),
    .io_addressOut_ready(queues_36_io_addressOut_ready),
    .io_addressOut_valid(queues_36_io_addressOut_valid),
    .io_addressOut_bits(queues_36_io_addressOut_bits)
  );
  contQueue_64 queues_37 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_37_clock),
    .reset(queues_37_reset),
    .io_addressIn_ready(queues_37_io_addressIn_ready),
    .io_addressIn_valid(queues_37_io_addressIn_valid),
    .io_addressIn_bits(queues_37_io_addressIn_bits),
    .io_addressOut_ready(queues_37_io_addressOut_ready),
    .io_addressOut_valid(queues_37_io_addressOut_valid),
    .io_addressOut_bits(queues_37_io_addressOut_bits)
  );
  contQueue_64 queues_38 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_38_clock),
    .reset(queues_38_reset),
    .io_addressIn_ready(queues_38_io_addressIn_ready),
    .io_addressIn_valid(queues_38_io_addressIn_valid),
    .io_addressIn_bits(queues_38_io_addressIn_bits),
    .io_addressOut_ready(queues_38_io_addressOut_ready),
    .io_addressOut_valid(queues_38_io_addressOut_valid),
    .io_addressOut_bits(queues_38_io_addressOut_bits)
  );
  contQueue_64 queues_39 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_39_clock),
    .reset(queues_39_reset),
    .io_addressIn_ready(queues_39_io_addressIn_ready),
    .io_addressIn_valid(queues_39_io_addressIn_valid),
    .io_addressIn_bits(queues_39_io_addressIn_bits),
    .io_addressOut_ready(queues_39_io_addressOut_ready),
    .io_addressOut_valid(queues_39_io_addressOut_valid),
    .io_addressOut_bits(queues_39_io_addressOut_bits)
  );
  contQueue_64 queues_40 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_40_clock),
    .reset(queues_40_reset),
    .io_addressIn_ready(queues_40_io_addressIn_ready),
    .io_addressIn_valid(queues_40_io_addressIn_valid),
    .io_addressIn_bits(queues_40_io_addressIn_bits),
    .io_addressOut_ready(queues_40_io_addressOut_ready),
    .io_addressOut_valid(queues_40_io_addressOut_valid),
    .io_addressOut_bits(queues_40_io_addressOut_bits)
  );
  contQueue_64 queues_41 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_41_clock),
    .reset(queues_41_reset),
    .io_addressIn_ready(queues_41_io_addressIn_ready),
    .io_addressIn_valid(queues_41_io_addressIn_valid),
    .io_addressIn_bits(queues_41_io_addressIn_bits),
    .io_addressOut_ready(queues_41_io_addressOut_ready),
    .io_addressOut_valid(queues_41_io_addressOut_valid),
    .io_addressOut_bits(queues_41_io_addressOut_bits)
  );
  contQueue_64 queues_42 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_42_clock),
    .reset(queues_42_reset),
    .io_addressIn_ready(queues_42_io_addressIn_ready),
    .io_addressIn_valid(queues_42_io_addressIn_valid),
    .io_addressIn_bits(queues_42_io_addressIn_bits),
    .io_addressOut_ready(queues_42_io_addressOut_ready),
    .io_addressOut_valid(queues_42_io_addressOut_valid),
    .io_addressOut_bits(queues_42_io_addressOut_bits)
  );
  contQueue_64 queues_43 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_43_clock),
    .reset(queues_43_reset),
    .io_addressIn_ready(queues_43_io_addressIn_ready),
    .io_addressIn_valid(queues_43_io_addressIn_valid),
    .io_addressIn_bits(queues_43_io_addressIn_bits),
    .io_addressOut_ready(queues_43_io_addressOut_ready),
    .io_addressOut_valid(queues_43_io_addressOut_valid),
    .io_addressOut_bits(queues_43_io_addressOut_bits)
  );
  contQueue_64 queues_44 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_44_clock),
    .reset(queues_44_reset),
    .io_addressIn_ready(queues_44_io_addressIn_ready),
    .io_addressIn_valid(queues_44_io_addressIn_valid),
    .io_addressIn_bits(queues_44_io_addressIn_bits),
    .io_addressOut_ready(queues_44_io_addressOut_ready),
    .io_addressOut_valid(queues_44_io_addressOut_valid),
    .io_addressOut_bits(queues_44_io_addressOut_bits)
  );
  contQueue_64 queues_45 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_45_clock),
    .reset(queues_45_reset),
    .io_addressIn_ready(queues_45_io_addressIn_ready),
    .io_addressIn_valid(queues_45_io_addressIn_valid),
    .io_addressIn_bits(queues_45_io_addressIn_bits),
    .io_addressOut_ready(queues_45_io_addressOut_ready),
    .io_addressOut_valid(queues_45_io_addressOut_valid),
    .io_addressOut_bits(queues_45_io_addressOut_bits)
  );
  contQueue_64 queues_46 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_46_clock),
    .reset(queues_46_reset),
    .io_addressIn_ready(queues_46_io_addressIn_ready),
    .io_addressIn_valid(queues_46_io_addressIn_valid),
    .io_addressIn_bits(queues_46_io_addressIn_bits),
    .io_addressOut_ready(queues_46_io_addressOut_ready),
    .io_addressOut_valid(queues_46_io_addressOut_valid),
    .io_addressOut_bits(queues_46_io_addressOut_bits)
  );
  contQueue_64 queues_47 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_47_clock),
    .reset(queues_47_reset),
    .io_addressIn_ready(queues_47_io_addressIn_ready),
    .io_addressIn_valid(queues_47_io_addressIn_valid),
    .io_addressIn_bits(queues_47_io_addressIn_bits),
    .io_addressOut_ready(queues_47_io_addressOut_ready),
    .io_addressOut_valid(queues_47_io_addressOut_valid),
    .io_addressOut_bits(queues_47_io_addressOut_bits)
  );
  contQueue_64 queues_48 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_48_clock),
    .reset(queues_48_reset),
    .io_addressIn_ready(queues_48_io_addressIn_ready),
    .io_addressIn_valid(queues_48_io_addressIn_valid),
    .io_addressIn_bits(queues_48_io_addressIn_bits),
    .io_addressOut_ready(queues_48_io_addressOut_ready),
    .io_addressOut_valid(queues_48_io_addressOut_valid),
    .io_addressOut_bits(queues_48_io_addressOut_bits)
  );
  contQueue_64 queues_49 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_49_clock),
    .reset(queues_49_reset),
    .io_addressIn_ready(queues_49_io_addressIn_ready),
    .io_addressIn_valid(queues_49_io_addressIn_valid),
    .io_addressIn_bits(queues_49_io_addressIn_bits),
    .io_addressOut_ready(queues_49_io_addressOut_ready),
    .io_addressOut_valid(queues_49_io_addressOut_valid),
    .io_addressOut_bits(queues_49_io_addressOut_bits)
  );
  contQueue_64 queues_50 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_50_clock),
    .reset(queues_50_reset),
    .io_addressIn_ready(queues_50_io_addressIn_ready),
    .io_addressIn_valid(queues_50_io_addressIn_valid),
    .io_addressIn_bits(queues_50_io_addressIn_bits),
    .io_addressOut_ready(queues_50_io_addressOut_ready),
    .io_addressOut_valid(queues_50_io_addressOut_valid),
    .io_addressOut_bits(queues_50_io_addressOut_bits)
  );
  contQueue_64 queues_51 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_51_clock),
    .reset(queues_51_reset),
    .io_addressIn_ready(queues_51_io_addressIn_ready),
    .io_addressIn_valid(queues_51_io_addressIn_valid),
    .io_addressIn_bits(queues_51_io_addressIn_bits),
    .io_addressOut_ready(queues_51_io_addressOut_ready),
    .io_addressOut_valid(queues_51_io_addressOut_valid),
    .io_addressOut_bits(queues_51_io_addressOut_bits)
  );
  contQueue_64 queues_52 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_52_clock),
    .reset(queues_52_reset),
    .io_addressIn_ready(queues_52_io_addressIn_ready),
    .io_addressIn_valid(queues_52_io_addressIn_valid),
    .io_addressIn_bits(queues_52_io_addressIn_bits),
    .io_addressOut_ready(queues_52_io_addressOut_ready),
    .io_addressOut_valid(queues_52_io_addressOut_valid),
    .io_addressOut_bits(queues_52_io_addressOut_bits)
  );
  contQueue_64 queues_53 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_53_clock),
    .reset(queues_53_reset),
    .io_addressIn_ready(queues_53_io_addressIn_ready),
    .io_addressIn_valid(queues_53_io_addressIn_valid),
    .io_addressIn_bits(queues_53_io_addressIn_bits),
    .io_addressOut_ready(queues_53_io_addressOut_ready),
    .io_addressOut_valid(queues_53_io_addressOut_valid),
    .io_addressOut_bits(queues_53_io_addressOut_bits)
  );
  contQueue_64 queues_54 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_54_clock),
    .reset(queues_54_reset),
    .io_addressIn_ready(queues_54_io_addressIn_ready),
    .io_addressIn_valid(queues_54_io_addressIn_valid),
    .io_addressIn_bits(queues_54_io_addressIn_bits),
    .io_addressOut_ready(queues_54_io_addressOut_ready),
    .io_addressOut_valid(queues_54_io_addressOut_valid),
    .io_addressOut_bits(queues_54_io_addressOut_bits)
  );
  contQueue_64 queues_55 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_55_clock),
    .reset(queues_55_reset),
    .io_addressIn_ready(queues_55_io_addressIn_ready),
    .io_addressIn_valid(queues_55_io_addressIn_valid),
    .io_addressIn_bits(queues_55_io_addressIn_bits),
    .io_addressOut_ready(queues_55_io_addressOut_ready),
    .io_addressOut_valid(queues_55_io_addressOut_valid),
    .io_addressOut_bits(queues_55_io_addressOut_bits)
  );
  contQueue_64 queues_56 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_56_clock),
    .reset(queues_56_reset),
    .io_addressIn_ready(queues_56_io_addressIn_ready),
    .io_addressIn_valid(queues_56_io_addressIn_valid),
    .io_addressIn_bits(queues_56_io_addressIn_bits),
    .io_addressOut_ready(queues_56_io_addressOut_ready),
    .io_addressOut_valid(queues_56_io_addressOut_valid),
    .io_addressOut_bits(queues_56_io_addressOut_bits)
  );
  contQueue_64 queues_57 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_57_clock),
    .reset(queues_57_reset),
    .io_addressIn_ready(queues_57_io_addressIn_ready),
    .io_addressIn_valid(queues_57_io_addressIn_valid),
    .io_addressIn_bits(queues_57_io_addressIn_bits),
    .io_addressOut_ready(queues_57_io_addressOut_ready),
    .io_addressOut_valid(queues_57_io_addressOut_valid),
    .io_addressOut_bits(queues_57_io_addressOut_bits)
  );
  contQueue_64 queues_58 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_58_clock),
    .reset(queues_58_reset),
    .io_addressIn_ready(queues_58_io_addressIn_ready),
    .io_addressIn_valid(queues_58_io_addressIn_valid),
    .io_addressIn_bits(queues_58_io_addressIn_bits),
    .io_addressOut_ready(queues_58_io_addressOut_ready),
    .io_addressOut_valid(queues_58_io_addressOut_valid),
    .io_addressOut_bits(queues_58_io_addressOut_bits)
  );
  contQueue_64 queues_59 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_59_clock),
    .reset(queues_59_reset),
    .io_addressIn_ready(queues_59_io_addressIn_ready),
    .io_addressIn_valid(queues_59_io_addressIn_valid),
    .io_addressIn_bits(queues_59_io_addressIn_bits),
    .io_addressOut_ready(queues_59_io_addressOut_ready),
    .io_addressOut_valid(queues_59_io_addressOut_valid),
    .io_addressOut_bits(queues_59_io_addressOut_bits)
  );
  contQueue_64 queues_60 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_60_clock),
    .reset(queues_60_reset),
    .io_addressIn_ready(queues_60_io_addressIn_ready),
    .io_addressIn_valid(queues_60_io_addressIn_valid),
    .io_addressIn_bits(queues_60_io_addressIn_bits),
    .io_addressOut_ready(queues_60_io_addressOut_ready),
    .io_addressOut_valid(queues_60_io_addressOut_valid),
    .io_addressOut_bits(queues_60_io_addressOut_bits)
  );
  contQueue_64 queues_61 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_61_clock),
    .reset(queues_61_reset),
    .io_addressIn_ready(queues_61_io_addressIn_ready),
    .io_addressIn_valid(queues_61_io_addressIn_valid),
    .io_addressIn_bits(queues_61_io_addressIn_bits),
    .io_addressOut_ready(queues_61_io_addressOut_ready),
    .io_addressOut_valid(queues_61_io_addressOut_valid),
    .io_addressOut_bits(queues_61_io_addressOut_bits)
  );
  contQueue_64 queues_62 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_62_clock),
    .reset(queues_62_reset),
    .io_addressIn_ready(queues_62_io_addressIn_ready),
    .io_addressIn_valid(queues_62_io_addressIn_valid),
    .io_addressIn_bits(queues_62_io_addressIn_bits),
    .io_addressOut_ready(queues_62_io_addressOut_ready),
    .io_addressOut_valid(queues_62_io_addressOut_valid),
    .io_addressOut_bits(queues_62_io_addressOut_bits)
  );
  contQueue_64 queues_63 ( // @[argRouteNetwork.scala 79:49]
    .clock(queues_63_clock),
    .reset(queues_63_reset),
    .io_addressIn_ready(queues_63_io_addressIn_ready),
    .io_addressIn_valid(queues_63_io_addressIn_valid),
    .io_addressIn_bits(queues_63_io_addressIn_bits),
    .io_addressOut_ready(queues_63_io_addressOut_ready),
    .io_addressOut_valid(queues_63_io_addressOut_valid),
    .io_addressOut_bits(queues_63_io_addressOut_bits)
  );
  assign io_connVAS_0_valid = virtNetworkUnits_0_io_vasAddressOut_valid; // @[argRouteNetwork.scala 107:46]
  assign io_connVAS_0_bits = virtNetworkUnits_0_io_vasAddressOut_bits; // @[argRouteNetwork.scala 107:46]
  assign io_connVAS_1_valid = virtNetworkUnits_1_io_vasAddressOut_valid; // @[argRouteNetwork.scala 107:46]
  assign io_connVAS_1_bits = virtNetworkUnits_1_io_vasAddressOut_bits; // @[argRouteNetwork.scala 107:46]
  assign io_connPE_0_ready = queues_0_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_1_ready = queues_1_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_2_ready = queues_2_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_3_ready = queues_3_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_4_ready = queues_4_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_5_ready = queues_5_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_6_ready = queues_6_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_7_ready = queues_7_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_8_ready = queues_8_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_9_ready = queues_9_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_10_ready = queues_10_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_11_ready = queues_11_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_12_ready = queues_12_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_13_ready = queues_13_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_14_ready = queues_14_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_15_ready = queues_15_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_16_ready = queues_16_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_17_ready = queues_17_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_18_ready = queues_18_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_19_ready = queues_19_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_20_ready = queues_20_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_21_ready = queues_21_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_22_ready = queues_22_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_23_ready = queues_23_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_24_ready = queues_24_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_25_ready = queues_25_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_26_ready = queues_26_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_27_ready = queues_27_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_28_ready = queues_28_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_29_ready = queues_29_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_30_ready = queues_30_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_31_ready = queues_31_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_32_ready = queues_32_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_33_ready = queues_33_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_34_ready = queues_34_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_35_ready = queues_35_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_36_ready = queues_36_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_37_ready = queues_37_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_38_ready = queues_38_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_39_ready = queues_39_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_40_ready = queues_40_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_41_ready = queues_41_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_42_ready = queues_42_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_43_ready = queues_43_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_44_ready = queues_44_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_45_ready = queues_45_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_46_ready = queues_46_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_47_ready = queues_47_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_48_ready = queues_48_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_49_ready = queues_49_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_50_ready = queues_50_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_51_ready = queues_51_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_52_ready = queues_52_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_53_ready = queues_53_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_54_ready = queues_54_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_55_ready = queues_55_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_56_ready = queues_56_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_57_ready = queues_57_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_58_ready = queues_58_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_59_ready = queues_59_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_60_ready = queues_60_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_61_ready = queues_61_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_62_ready = queues_62_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign io_connPE_63_ready = queues_63_io_addressIn_ready; // @[argRouteNetwork.scala 83:21]
  assign networkUnits_0_clock = clock;
  assign networkUnits_0_reset = reset;
  assign networkUnits_0_io_addressIn_valid = networkUnits_1_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_0_io_addressIn_bits = networkUnits_1_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_0_io_peAddress_valid = queues_0_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_0_io_peAddress_bits = queues_0_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_0_io_addressOut_ready = virtNetworkUnits_1_io_addressIn_ready; // @[argRouteNetwork.scala 99:47]
  assign networkUnits_1_clock = clock;
  assign networkUnits_1_reset = reset;
  assign networkUnits_1_io_addressIn_valid = networkUnits_2_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_1_io_addressIn_bits = networkUnits_2_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_1_io_peAddress_valid = queues_1_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_1_io_peAddress_bits = queues_1_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_1_io_addressOut_ready = networkUnits_0_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_2_clock = clock;
  assign networkUnits_2_reset = reset;
  assign networkUnits_2_io_addressIn_valid = networkUnits_3_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_2_io_addressIn_bits = networkUnits_3_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_2_io_peAddress_valid = queues_2_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_2_io_peAddress_bits = queues_2_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_2_io_addressOut_ready = networkUnits_1_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_3_clock = clock;
  assign networkUnits_3_reset = reset;
  assign networkUnits_3_io_addressIn_valid = networkUnits_4_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_3_io_addressIn_bits = networkUnits_4_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_3_io_peAddress_valid = queues_3_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_3_io_peAddress_bits = queues_3_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_3_io_addressOut_ready = networkUnits_2_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_4_clock = clock;
  assign networkUnits_4_reset = reset;
  assign networkUnits_4_io_addressIn_valid = networkUnits_5_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_4_io_addressIn_bits = networkUnits_5_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_4_io_peAddress_valid = queues_4_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_4_io_peAddress_bits = queues_4_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_4_io_addressOut_ready = networkUnits_3_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_5_clock = clock;
  assign networkUnits_5_reset = reset;
  assign networkUnits_5_io_addressIn_valid = networkUnits_6_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_5_io_addressIn_bits = networkUnits_6_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_5_io_peAddress_valid = queues_5_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_5_io_peAddress_bits = queues_5_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_5_io_addressOut_ready = networkUnits_4_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_6_clock = clock;
  assign networkUnits_6_reset = reset;
  assign networkUnits_6_io_addressIn_valid = networkUnits_7_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_6_io_addressIn_bits = networkUnits_7_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_6_io_peAddress_valid = queues_6_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_6_io_peAddress_bits = queues_6_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_6_io_addressOut_ready = networkUnits_5_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_7_clock = clock;
  assign networkUnits_7_reset = reset;
  assign networkUnits_7_io_addressIn_valid = networkUnits_8_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_7_io_addressIn_bits = networkUnits_8_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_7_io_peAddress_valid = queues_7_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_7_io_peAddress_bits = queues_7_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_7_io_addressOut_ready = networkUnits_6_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_8_clock = clock;
  assign networkUnits_8_reset = reset;
  assign networkUnits_8_io_addressIn_valid = networkUnits_9_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_8_io_addressIn_bits = networkUnits_9_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_8_io_peAddress_valid = queues_8_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_8_io_peAddress_bits = queues_8_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_8_io_addressOut_ready = networkUnits_7_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_9_clock = clock;
  assign networkUnits_9_reset = reset;
  assign networkUnits_9_io_addressIn_valid = networkUnits_10_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_9_io_addressIn_bits = networkUnits_10_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_9_io_peAddress_valid = queues_9_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_9_io_peAddress_bits = queues_9_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_9_io_addressOut_ready = networkUnits_8_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_10_clock = clock;
  assign networkUnits_10_reset = reset;
  assign networkUnits_10_io_addressIn_valid = networkUnits_11_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_10_io_addressIn_bits = networkUnits_11_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_10_io_peAddress_valid = queues_10_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_10_io_peAddress_bits = queues_10_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_10_io_addressOut_ready = networkUnits_9_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_11_clock = clock;
  assign networkUnits_11_reset = reset;
  assign networkUnits_11_io_addressIn_valid = networkUnits_12_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_11_io_addressIn_bits = networkUnits_12_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_11_io_peAddress_valid = queues_11_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_11_io_peAddress_bits = queues_11_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_11_io_addressOut_ready = networkUnits_10_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_12_clock = clock;
  assign networkUnits_12_reset = reset;
  assign networkUnits_12_io_addressIn_valid = networkUnits_13_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_12_io_addressIn_bits = networkUnits_13_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_12_io_peAddress_valid = queues_12_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_12_io_peAddress_bits = queues_12_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_12_io_addressOut_ready = networkUnits_11_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_13_clock = clock;
  assign networkUnits_13_reset = reset;
  assign networkUnits_13_io_addressIn_valid = networkUnits_14_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_13_io_addressIn_bits = networkUnits_14_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_13_io_peAddress_valid = queues_13_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_13_io_peAddress_bits = queues_13_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_13_io_addressOut_ready = networkUnits_12_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_14_clock = clock;
  assign networkUnits_14_reset = reset;
  assign networkUnits_14_io_addressIn_valid = networkUnits_15_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_14_io_addressIn_bits = networkUnits_15_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_14_io_peAddress_valid = queues_14_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_14_io_peAddress_bits = queues_14_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_14_io_addressOut_ready = networkUnits_13_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_15_clock = clock;
  assign networkUnits_15_reset = reset;
  assign networkUnits_15_io_addressIn_valid = networkUnits_16_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_15_io_addressIn_bits = networkUnits_16_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_15_io_peAddress_valid = queues_15_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_15_io_peAddress_bits = queues_15_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_15_io_addressOut_ready = networkUnits_14_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_16_clock = clock;
  assign networkUnits_16_reset = reset;
  assign networkUnits_16_io_addressIn_valid = networkUnits_17_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_16_io_addressIn_bits = networkUnits_17_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_16_io_peAddress_valid = queues_16_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_16_io_peAddress_bits = queues_16_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_16_io_addressOut_ready = networkUnits_15_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_17_clock = clock;
  assign networkUnits_17_reset = reset;
  assign networkUnits_17_io_addressIn_valid = networkUnits_18_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_17_io_addressIn_bits = networkUnits_18_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_17_io_peAddress_valid = queues_17_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_17_io_peAddress_bits = queues_17_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_17_io_addressOut_ready = networkUnits_16_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_18_clock = clock;
  assign networkUnits_18_reset = reset;
  assign networkUnits_18_io_addressIn_valid = networkUnits_19_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_18_io_addressIn_bits = networkUnits_19_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_18_io_peAddress_valid = queues_18_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_18_io_peAddress_bits = queues_18_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_18_io_addressOut_ready = networkUnits_17_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_19_clock = clock;
  assign networkUnits_19_reset = reset;
  assign networkUnits_19_io_addressIn_valid = networkUnits_20_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_19_io_addressIn_bits = networkUnits_20_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_19_io_peAddress_valid = queues_19_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_19_io_peAddress_bits = queues_19_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_19_io_addressOut_ready = networkUnits_18_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_20_clock = clock;
  assign networkUnits_20_reset = reset;
  assign networkUnits_20_io_addressIn_valid = networkUnits_21_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_20_io_addressIn_bits = networkUnits_21_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_20_io_peAddress_valid = queues_20_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_20_io_peAddress_bits = queues_20_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_20_io_addressOut_ready = networkUnits_19_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_21_clock = clock;
  assign networkUnits_21_reset = reset;
  assign networkUnits_21_io_addressIn_valid = networkUnits_22_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_21_io_addressIn_bits = networkUnits_22_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_21_io_peAddress_valid = queues_21_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_21_io_peAddress_bits = queues_21_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_21_io_addressOut_ready = networkUnits_20_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_22_clock = clock;
  assign networkUnits_22_reset = reset;
  assign networkUnits_22_io_addressIn_valid = networkUnits_23_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_22_io_addressIn_bits = networkUnits_23_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_22_io_peAddress_valid = queues_22_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_22_io_peAddress_bits = queues_22_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_22_io_addressOut_ready = networkUnits_21_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_23_clock = clock;
  assign networkUnits_23_reset = reset;
  assign networkUnits_23_io_addressIn_valid = networkUnits_24_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_23_io_addressIn_bits = networkUnits_24_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_23_io_peAddress_valid = queues_23_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_23_io_peAddress_bits = queues_23_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_23_io_addressOut_ready = networkUnits_22_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_24_clock = clock;
  assign networkUnits_24_reset = reset;
  assign networkUnits_24_io_addressIn_valid = networkUnits_25_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_24_io_addressIn_bits = networkUnits_25_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_24_io_peAddress_valid = queues_24_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_24_io_peAddress_bits = queues_24_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_24_io_addressOut_ready = networkUnits_23_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_25_clock = clock;
  assign networkUnits_25_reset = reset;
  assign networkUnits_25_io_addressIn_valid = networkUnits_26_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_25_io_addressIn_bits = networkUnits_26_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_25_io_peAddress_valid = queues_25_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_25_io_peAddress_bits = queues_25_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_25_io_addressOut_ready = networkUnits_24_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_26_clock = clock;
  assign networkUnits_26_reset = reset;
  assign networkUnits_26_io_addressIn_valid = networkUnits_27_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_26_io_addressIn_bits = networkUnits_27_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_26_io_peAddress_valid = queues_26_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_26_io_peAddress_bits = queues_26_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_26_io_addressOut_ready = networkUnits_25_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_27_clock = clock;
  assign networkUnits_27_reset = reset;
  assign networkUnits_27_io_addressIn_valid = networkUnits_28_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_27_io_addressIn_bits = networkUnits_28_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_27_io_peAddress_valid = queues_27_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_27_io_peAddress_bits = queues_27_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_27_io_addressOut_ready = networkUnits_26_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_28_clock = clock;
  assign networkUnits_28_reset = reset;
  assign networkUnits_28_io_addressIn_valid = networkUnits_29_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_28_io_addressIn_bits = networkUnits_29_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_28_io_peAddress_valid = queues_28_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_28_io_peAddress_bits = queues_28_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_28_io_addressOut_ready = networkUnits_27_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_29_clock = clock;
  assign networkUnits_29_reset = reset;
  assign networkUnits_29_io_addressIn_valid = networkUnits_30_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_29_io_addressIn_bits = networkUnits_30_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_29_io_peAddress_valid = queues_29_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_29_io_peAddress_bits = queues_29_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_29_io_addressOut_ready = networkUnits_28_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_30_clock = clock;
  assign networkUnits_30_reset = reset;
  assign networkUnits_30_io_addressIn_valid = networkUnits_31_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_30_io_addressIn_bits = networkUnits_31_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_30_io_peAddress_valid = queues_30_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_30_io_peAddress_bits = queues_30_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_30_io_addressOut_ready = networkUnits_29_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_31_clock = clock;
  assign networkUnits_31_reset = reset;
  assign networkUnits_31_io_addressIn_valid = networkUnits_32_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_31_io_addressIn_bits = networkUnits_32_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_31_io_peAddress_valid = queues_31_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_31_io_peAddress_bits = queues_31_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_31_io_addressOut_ready = networkUnits_30_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_32_clock = clock;
  assign networkUnits_32_reset = reset;
  assign networkUnits_32_io_addressIn_valid = networkUnits_33_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_32_io_addressIn_bits = networkUnits_33_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_32_io_peAddress_valid = queues_32_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_32_io_peAddress_bits = queues_32_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_32_io_addressOut_ready = networkUnits_31_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_33_clock = clock;
  assign networkUnits_33_reset = reset;
  assign networkUnits_33_io_addressIn_valid = networkUnits_34_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_33_io_addressIn_bits = networkUnits_34_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_33_io_peAddress_valid = queues_33_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_33_io_peAddress_bits = queues_33_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_33_io_addressOut_ready = networkUnits_32_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_34_clock = clock;
  assign networkUnits_34_reset = reset;
  assign networkUnits_34_io_addressIn_valid = networkUnits_35_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_34_io_addressIn_bits = networkUnits_35_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_34_io_peAddress_valid = queues_34_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_34_io_peAddress_bits = queues_34_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_34_io_addressOut_ready = networkUnits_33_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_35_clock = clock;
  assign networkUnits_35_reset = reset;
  assign networkUnits_35_io_addressIn_valid = networkUnits_36_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_35_io_addressIn_bits = networkUnits_36_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_35_io_peAddress_valid = queues_35_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_35_io_peAddress_bits = queues_35_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_35_io_addressOut_ready = networkUnits_34_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_36_clock = clock;
  assign networkUnits_36_reset = reset;
  assign networkUnits_36_io_addressIn_valid = networkUnits_37_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_36_io_addressIn_bits = networkUnits_37_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_36_io_peAddress_valid = queues_36_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_36_io_peAddress_bits = queues_36_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_36_io_addressOut_ready = networkUnits_35_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_37_clock = clock;
  assign networkUnits_37_reset = reset;
  assign networkUnits_37_io_addressIn_valid = networkUnits_38_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_37_io_addressIn_bits = networkUnits_38_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_37_io_peAddress_valid = queues_37_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_37_io_peAddress_bits = queues_37_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_37_io_addressOut_ready = networkUnits_36_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_38_clock = clock;
  assign networkUnits_38_reset = reset;
  assign networkUnits_38_io_addressIn_valid = networkUnits_39_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_38_io_addressIn_bits = networkUnits_39_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_38_io_peAddress_valid = queues_38_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_38_io_peAddress_bits = queues_38_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_38_io_addressOut_ready = networkUnits_37_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_39_clock = clock;
  assign networkUnits_39_reset = reset;
  assign networkUnits_39_io_addressIn_valid = networkUnits_40_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_39_io_addressIn_bits = networkUnits_40_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_39_io_peAddress_valid = queues_39_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_39_io_peAddress_bits = queues_39_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_39_io_addressOut_ready = networkUnits_38_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_40_clock = clock;
  assign networkUnits_40_reset = reset;
  assign networkUnits_40_io_addressIn_valid = networkUnits_41_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_40_io_addressIn_bits = networkUnits_41_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_40_io_peAddress_valid = queues_40_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_40_io_peAddress_bits = queues_40_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_40_io_addressOut_ready = networkUnits_39_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_41_clock = clock;
  assign networkUnits_41_reset = reset;
  assign networkUnits_41_io_addressIn_valid = networkUnits_42_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_41_io_addressIn_bits = networkUnits_42_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_41_io_peAddress_valid = queues_41_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_41_io_peAddress_bits = queues_41_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_41_io_addressOut_ready = networkUnits_40_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_42_clock = clock;
  assign networkUnits_42_reset = reset;
  assign networkUnits_42_io_addressIn_valid = networkUnits_43_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_42_io_addressIn_bits = networkUnits_43_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_42_io_peAddress_valid = queues_42_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_42_io_peAddress_bits = queues_42_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_42_io_addressOut_ready = networkUnits_41_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_43_clock = clock;
  assign networkUnits_43_reset = reset;
  assign networkUnits_43_io_addressIn_valid = networkUnits_44_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_43_io_addressIn_bits = networkUnits_44_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_43_io_peAddress_valid = queues_43_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_43_io_peAddress_bits = queues_43_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_43_io_addressOut_ready = networkUnits_42_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_44_clock = clock;
  assign networkUnits_44_reset = reset;
  assign networkUnits_44_io_addressIn_valid = networkUnits_45_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_44_io_addressIn_bits = networkUnits_45_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_44_io_peAddress_valid = queues_44_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_44_io_peAddress_bits = queues_44_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_44_io_addressOut_ready = networkUnits_43_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_45_clock = clock;
  assign networkUnits_45_reset = reset;
  assign networkUnits_45_io_addressIn_valid = networkUnits_46_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_45_io_addressIn_bits = networkUnits_46_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_45_io_peAddress_valid = queues_45_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_45_io_peAddress_bits = queues_45_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_45_io_addressOut_ready = networkUnits_44_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_46_clock = clock;
  assign networkUnits_46_reset = reset;
  assign networkUnits_46_io_addressIn_valid = networkUnits_47_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_46_io_addressIn_bits = networkUnits_47_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_46_io_peAddress_valid = queues_46_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_46_io_peAddress_bits = queues_46_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_46_io_addressOut_ready = networkUnits_45_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_47_clock = clock;
  assign networkUnits_47_reset = reset;
  assign networkUnits_47_io_addressIn_valid = networkUnits_48_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_47_io_addressIn_bits = networkUnits_48_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_47_io_peAddress_valid = queues_47_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_47_io_peAddress_bits = queues_47_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_47_io_addressOut_ready = networkUnits_46_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_48_clock = clock;
  assign networkUnits_48_reset = reset;
  assign networkUnits_48_io_addressIn_valid = networkUnits_49_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_48_io_addressIn_bits = networkUnits_49_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_48_io_peAddress_valid = queues_48_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_48_io_peAddress_bits = queues_48_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_48_io_addressOut_ready = networkUnits_47_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_49_clock = clock;
  assign networkUnits_49_reset = reset;
  assign networkUnits_49_io_addressIn_valid = networkUnits_50_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_49_io_addressIn_bits = networkUnits_50_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_49_io_peAddress_valid = queues_49_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_49_io_peAddress_bits = queues_49_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_49_io_addressOut_ready = networkUnits_48_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_50_clock = clock;
  assign networkUnits_50_reset = reset;
  assign networkUnits_50_io_addressIn_valid = networkUnits_51_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_50_io_addressIn_bits = networkUnits_51_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_50_io_peAddress_valid = queues_50_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_50_io_peAddress_bits = queues_50_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_50_io_addressOut_ready = networkUnits_49_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_51_clock = clock;
  assign networkUnits_51_reset = reset;
  assign networkUnits_51_io_addressIn_valid = networkUnits_52_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_51_io_addressIn_bits = networkUnits_52_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_51_io_peAddress_valid = queues_51_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_51_io_peAddress_bits = queues_51_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_51_io_addressOut_ready = networkUnits_50_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_52_clock = clock;
  assign networkUnits_52_reset = reset;
  assign networkUnits_52_io_addressIn_valid = networkUnits_53_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_52_io_addressIn_bits = networkUnits_53_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_52_io_peAddress_valid = queues_52_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_52_io_peAddress_bits = queues_52_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_52_io_addressOut_ready = networkUnits_51_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_53_clock = clock;
  assign networkUnits_53_reset = reset;
  assign networkUnits_53_io_addressIn_valid = networkUnits_54_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_53_io_addressIn_bits = networkUnits_54_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_53_io_peAddress_valid = queues_53_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_53_io_peAddress_bits = queues_53_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_53_io_addressOut_ready = networkUnits_52_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_54_clock = clock;
  assign networkUnits_54_reset = reset;
  assign networkUnits_54_io_addressIn_valid = networkUnits_55_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_54_io_addressIn_bits = networkUnits_55_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_54_io_peAddress_valid = queues_54_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_54_io_peAddress_bits = queues_54_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_54_io_addressOut_ready = networkUnits_53_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_55_clock = clock;
  assign networkUnits_55_reset = reset;
  assign networkUnits_55_io_addressIn_valid = networkUnits_56_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_55_io_addressIn_bits = networkUnits_56_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_55_io_peAddress_valid = queues_55_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_55_io_peAddress_bits = queues_55_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_55_io_addressOut_ready = networkUnits_54_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_56_clock = clock;
  assign networkUnits_56_reset = reset;
  assign networkUnits_56_io_addressIn_valid = networkUnits_57_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_56_io_addressIn_bits = networkUnits_57_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_56_io_peAddress_valid = queues_56_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_56_io_peAddress_bits = queues_56_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_56_io_addressOut_ready = networkUnits_55_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_57_clock = clock;
  assign networkUnits_57_reset = reset;
  assign networkUnits_57_io_addressIn_valid = networkUnits_58_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_57_io_addressIn_bits = networkUnits_58_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_57_io_peAddress_valid = queues_57_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_57_io_peAddress_bits = queues_57_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_57_io_addressOut_ready = networkUnits_56_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_58_clock = clock;
  assign networkUnits_58_reset = reset;
  assign networkUnits_58_io_addressIn_valid = networkUnits_59_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_58_io_addressIn_bits = networkUnits_59_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_58_io_peAddress_valid = queues_58_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_58_io_peAddress_bits = queues_58_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_58_io_addressOut_ready = networkUnits_57_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_59_clock = clock;
  assign networkUnits_59_reset = reset;
  assign networkUnits_59_io_addressIn_valid = networkUnits_60_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_59_io_addressIn_bits = networkUnits_60_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_59_io_peAddress_valid = queues_59_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_59_io_peAddress_bits = queues_59_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_59_io_addressOut_ready = networkUnits_58_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_60_clock = clock;
  assign networkUnits_60_reset = reset;
  assign networkUnits_60_io_addressIn_valid = networkUnits_61_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_60_io_addressIn_bits = networkUnits_61_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_60_io_peAddress_valid = queues_60_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_60_io_peAddress_bits = queues_60_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_60_io_addressOut_ready = networkUnits_59_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_61_clock = clock;
  assign networkUnits_61_reset = reset;
  assign networkUnits_61_io_addressIn_valid = networkUnits_62_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_61_io_addressIn_bits = networkUnits_62_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_61_io_peAddress_valid = queues_61_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_61_io_peAddress_bits = queues_61_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_61_io_addressOut_ready = networkUnits_60_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_62_clock = clock;
  assign networkUnits_62_reset = reset;
  assign networkUnits_62_io_addressIn_valid = networkUnits_63_io_addressOut_valid; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_62_io_addressIn_bits = networkUnits_63_io_addressOut_bits; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_62_io_peAddress_valid = queues_62_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_62_io_peAddress_bits = queues_62_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_62_io_addressOut_ready = networkUnits_61_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign networkUnits_63_clock = clock;
  assign networkUnits_63_reset = reset;
  assign networkUnits_63_io_addressIn_valid = 1'h0; // @[argRouteNetwork.scala 95:50]
  assign networkUnits_63_io_addressIn_bits = 64'h0; // @[argRouteNetwork.scala 42:{46,46}]
  assign networkUnits_63_io_peAddress_valid = queues_63_io_addressOut_valid; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_63_io_peAddress_bits = queues_63_io_addressOut_bits; // @[argRouteNetwork.scala 92:38]
  assign networkUnits_63_io_addressOut_ready = networkUnits_62_io_addressIn_ready; // @[argRouteNetwork.scala 88:38]
  assign virtNetworkUnits_0_clock = clock;
  assign virtNetworkUnits_0_reset = reset;
  assign virtNetworkUnits_0_io_addressIn_valid = virtNetworkUnits_1_io_addressOut_valid; // @[argRouteNetwork.scala 103:42]
  assign virtNetworkUnits_0_io_addressIn_bits = virtNetworkUnits_1_io_addressOut_bits; // @[argRouteNetwork.scala 103:42]
  assign virtNetworkUnits_0_io_vasAddressOut_ready = io_connVAS_0_ready; // @[argRouteNetwork.scala 107:46]
  assign virtNetworkUnits_1_clock = clock;
  assign virtNetworkUnits_1_reset = reset;
  assign virtNetworkUnits_1_io_addressIn_valid = networkUnits_0_io_addressOut_valid; // @[argRouteNetwork.scala 99:47]
  assign virtNetworkUnits_1_io_addressIn_bits = networkUnits_0_io_addressOut_bits; // @[argRouteNetwork.scala 99:47]
  assign virtNetworkUnits_1_io_vasAddressOut_ready = io_connVAS_1_ready; // @[argRouteNetwork.scala 107:46]
  assign virtNetworkUnits_1_io_addressOut_ready = virtNetworkUnits_0_io_addressIn_ready; // @[argRouteNetwork.scala 103:42]
  assign queues_0_clock = clock;
  assign queues_0_reset = reset;
  assign queues_0_io_addressIn_valid = io_connPE_0_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_0_io_addressIn_bits = io_connPE_0_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_0_io_addressOut_ready = networkUnits_0_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_1_clock = clock;
  assign queues_1_reset = reset;
  assign queues_1_io_addressIn_valid = io_connPE_1_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_1_io_addressIn_bits = io_connPE_1_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_1_io_addressOut_ready = networkUnits_1_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_2_clock = clock;
  assign queues_2_reset = reset;
  assign queues_2_io_addressIn_valid = io_connPE_2_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_2_io_addressIn_bits = io_connPE_2_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_2_io_addressOut_ready = networkUnits_2_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_3_clock = clock;
  assign queues_3_reset = reset;
  assign queues_3_io_addressIn_valid = io_connPE_3_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_3_io_addressIn_bits = io_connPE_3_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_3_io_addressOut_ready = networkUnits_3_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_4_clock = clock;
  assign queues_4_reset = reset;
  assign queues_4_io_addressIn_valid = io_connPE_4_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_4_io_addressIn_bits = io_connPE_4_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_4_io_addressOut_ready = networkUnits_4_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_5_clock = clock;
  assign queues_5_reset = reset;
  assign queues_5_io_addressIn_valid = io_connPE_5_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_5_io_addressIn_bits = io_connPE_5_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_5_io_addressOut_ready = networkUnits_5_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_6_clock = clock;
  assign queues_6_reset = reset;
  assign queues_6_io_addressIn_valid = io_connPE_6_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_6_io_addressIn_bits = io_connPE_6_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_6_io_addressOut_ready = networkUnits_6_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_7_clock = clock;
  assign queues_7_reset = reset;
  assign queues_7_io_addressIn_valid = io_connPE_7_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_7_io_addressIn_bits = io_connPE_7_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_7_io_addressOut_ready = networkUnits_7_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_8_clock = clock;
  assign queues_8_reset = reset;
  assign queues_8_io_addressIn_valid = io_connPE_8_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_8_io_addressIn_bits = io_connPE_8_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_8_io_addressOut_ready = networkUnits_8_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_9_clock = clock;
  assign queues_9_reset = reset;
  assign queues_9_io_addressIn_valid = io_connPE_9_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_9_io_addressIn_bits = io_connPE_9_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_9_io_addressOut_ready = networkUnits_9_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_10_clock = clock;
  assign queues_10_reset = reset;
  assign queues_10_io_addressIn_valid = io_connPE_10_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_10_io_addressIn_bits = io_connPE_10_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_10_io_addressOut_ready = networkUnits_10_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_11_clock = clock;
  assign queues_11_reset = reset;
  assign queues_11_io_addressIn_valid = io_connPE_11_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_11_io_addressIn_bits = io_connPE_11_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_11_io_addressOut_ready = networkUnits_11_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_12_clock = clock;
  assign queues_12_reset = reset;
  assign queues_12_io_addressIn_valid = io_connPE_12_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_12_io_addressIn_bits = io_connPE_12_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_12_io_addressOut_ready = networkUnits_12_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_13_clock = clock;
  assign queues_13_reset = reset;
  assign queues_13_io_addressIn_valid = io_connPE_13_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_13_io_addressIn_bits = io_connPE_13_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_13_io_addressOut_ready = networkUnits_13_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_14_clock = clock;
  assign queues_14_reset = reset;
  assign queues_14_io_addressIn_valid = io_connPE_14_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_14_io_addressIn_bits = io_connPE_14_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_14_io_addressOut_ready = networkUnits_14_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_15_clock = clock;
  assign queues_15_reset = reset;
  assign queues_15_io_addressIn_valid = io_connPE_15_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_15_io_addressIn_bits = io_connPE_15_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_15_io_addressOut_ready = networkUnits_15_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_16_clock = clock;
  assign queues_16_reset = reset;
  assign queues_16_io_addressIn_valid = io_connPE_16_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_16_io_addressIn_bits = io_connPE_16_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_16_io_addressOut_ready = networkUnits_16_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_17_clock = clock;
  assign queues_17_reset = reset;
  assign queues_17_io_addressIn_valid = io_connPE_17_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_17_io_addressIn_bits = io_connPE_17_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_17_io_addressOut_ready = networkUnits_17_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_18_clock = clock;
  assign queues_18_reset = reset;
  assign queues_18_io_addressIn_valid = io_connPE_18_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_18_io_addressIn_bits = io_connPE_18_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_18_io_addressOut_ready = networkUnits_18_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_19_clock = clock;
  assign queues_19_reset = reset;
  assign queues_19_io_addressIn_valid = io_connPE_19_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_19_io_addressIn_bits = io_connPE_19_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_19_io_addressOut_ready = networkUnits_19_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_20_clock = clock;
  assign queues_20_reset = reset;
  assign queues_20_io_addressIn_valid = io_connPE_20_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_20_io_addressIn_bits = io_connPE_20_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_20_io_addressOut_ready = networkUnits_20_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_21_clock = clock;
  assign queues_21_reset = reset;
  assign queues_21_io_addressIn_valid = io_connPE_21_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_21_io_addressIn_bits = io_connPE_21_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_21_io_addressOut_ready = networkUnits_21_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_22_clock = clock;
  assign queues_22_reset = reset;
  assign queues_22_io_addressIn_valid = io_connPE_22_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_22_io_addressIn_bits = io_connPE_22_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_22_io_addressOut_ready = networkUnits_22_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_23_clock = clock;
  assign queues_23_reset = reset;
  assign queues_23_io_addressIn_valid = io_connPE_23_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_23_io_addressIn_bits = io_connPE_23_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_23_io_addressOut_ready = networkUnits_23_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_24_clock = clock;
  assign queues_24_reset = reset;
  assign queues_24_io_addressIn_valid = io_connPE_24_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_24_io_addressIn_bits = io_connPE_24_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_24_io_addressOut_ready = networkUnits_24_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_25_clock = clock;
  assign queues_25_reset = reset;
  assign queues_25_io_addressIn_valid = io_connPE_25_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_25_io_addressIn_bits = io_connPE_25_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_25_io_addressOut_ready = networkUnits_25_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_26_clock = clock;
  assign queues_26_reset = reset;
  assign queues_26_io_addressIn_valid = io_connPE_26_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_26_io_addressIn_bits = io_connPE_26_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_26_io_addressOut_ready = networkUnits_26_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_27_clock = clock;
  assign queues_27_reset = reset;
  assign queues_27_io_addressIn_valid = io_connPE_27_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_27_io_addressIn_bits = io_connPE_27_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_27_io_addressOut_ready = networkUnits_27_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_28_clock = clock;
  assign queues_28_reset = reset;
  assign queues_28_io_addressIn_valid = io_connPE_28_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_28_io_addressIn_bits = io_connPE_28_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_28_io_addressOut_ready = networkUnits_28_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_29_clock = clock;
  assign queues_29_reset = reset;
  assign queues_29_io_addressIn_valid = io_connPE_29_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_29_io_addressIn_bits = io_connPE_29_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_29_io_addressOut_ready = networkUnits_29_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_30_clock = clock;
  assign queues_30_reset = reset;
  assign queues_30_io_addressIn_valid = io_connPE_30_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_30_io_addressIn_bits = io_connPE_30_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_30_io_addressOut_ready = networkUnits_30_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_31_clock = clock;
  assign queues_31_reset = reset;
  assign queues_31_io_addressIn_valid = io_connPE_31_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_31_io_addressIn_bits = io_connPE_31_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_31_io_addressOut_ready = networkUnits_31_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_32_clock = clock;
  assign queues_32_reset = reset;
  assign queues_32_io_addressIn_valid = io_connPE_32_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_32_io_addressIn_bits = io_connPE_32_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_32_io_addressOut_ready = networkUnits_32_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_33_clock = clock;
  assign queues_33_reset = reset;
  assign queues_33_io_addressIn_valid = io_connPE_33_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_33_io_addressIn_bits = io_connPE_33_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_33_io_addressOut_ready = networkUnits_33_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_34_clock = clock;
  assign queues_34_reset = reset;
  assign queues_34_io_addressIn_valid = io_connPE_34_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_34_io_addressIn_bits = io_connPE_34_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_34_io_addressOut_ready = networkUnits_34_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_35_clock = clock;
  assign queues_35_reset = reset;
  assign queues_35_io_addressIn_valid = io_connPE_35_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_35_io_addressIn_bits = io_connPE_35_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_35_io_addressOut_ready = networkUnits_35_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_36_clock = clock;
  assign queues_36_reset = reset;
  assign queues_36_io_addressIn_valid = io_connPE_36_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_36_io_addressIn_bits = io_connPE_36_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_36_io_addressOut_ready = networkUnits_36_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_37_clock = clock;
  assign queues_37_reset = reset;
  assign queues_37_io_addressIn_valid = io_connPE_37_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_37_io_addressIn_bits = io_connPE_37_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_37_io_addressOut_ready = networkUnits_37_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_38_clock = clock;
  assign queues_38_reset = reset;
  assign queues_38_io_addressIn_valid = io_connPE_38_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_38_io_addressIn_bits = io_connPE_38_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_38_io_addressOut_ready = networkUnits_38_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_39_clock = clock;
  assign queues_39_reset = reset;
  assign queues_39_io_addressIn_valid = io_connPE_39_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_39_io_addressIn_bits = io_connPE_39_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_39_io_addressOut_ready = networkUnits_39_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_40_clock = clock;
  assign queues_40_reset = reset;
  assign queues_40_io_addressIn_valid = io_connPE_40_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_40_io_addressIn_bits = io_connPE_40_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_40_io_addressOut_ready = networkUnits_40_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_41_clock = clock;
  assign queues_41_reset = reset;
  assign queues_41_io_addressIn_valid = io_connPE_41_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_41_io_addressIn_bits = io_connPE_41_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_41_io_addressOut_ready = networkUnits_41_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_42_clock = clock;
  assign queues_42_reset = reset;
  assign queues_42_io_addressIn_valid = io_connPE_42_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_42_io_addressIn_bits = io_connPE_42_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_42_io_addressOut_ready = networkUnits_42_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_43_clock = clock;
  assign queues_43_reset = reset;
  assign queues_43_io_addressIn_valid = io_connPE_43_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_43_io_addressIn_bits = io_connPE_43_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_43_io_addressOut_ready = networkUnits_43_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_44_clock = clock;
  assign queues_44_reset = reset;
  assign queues_44_io_addressIn_valid = io_connPE_44_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_44_io_addressIn_bits = io_connPE_44_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_44_io_addressOut_ready = networkUnits_44_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_45_clock = clock;
  assign queues_45_reset = reset;
  assign queues_45_io_addressIn_valid = io_connPE_45_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_45_io_addressIn_bits = io_connPE_45_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_45_io_addressOut_ready = networkUnits_45_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_46_clock = clock;
  assign queues_46_reset = reset;
  assign queues_46_io_addressIn_valid = io_connPE_46_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_46_io_addressIn_bits = io_connPE_46_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_46_io_addressOut_ready = networkUnits_46_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_47_clock = clock;
  assign queues_47_reset = reset;
  assign queues_47_io_addressIn_valid = io_connPE_47_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_47_io_addressIn_bits = io_connPE_47_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_47_io_addressOut_ready = networkUnits_47_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_48_clock = clock;
  assign queues_48_reset = reset;
  assign queues_48_io_addressIn_valid = io_connPE_48_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_48_io_addressIn_bits = io_connPE_48_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_48_io_addressOut_ready = networkUnits_48_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_49_clock = clock;
  assign queues_49_reset = reset;
  assign queues_49_io_addressIn_valid = io_connPE_49_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_49_io_addressIn_bits = io_connPE_49_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_49_io_addressOut_ready = networkUnits_49_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_50_clock = clock;
  assign queues_50_reset = reset;
  assign queues_50_io_addressIn_valid = io_connPE_50_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_50_io_addressIn_bits = io_connPE_50_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_50_io_addressOut_ready = networkUnits_50_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_51_clock = clock;
  assign queues_51_reset = reset;
  assign queues_51_io_addressIn_valid = io_connPE_51_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_51_io_addressIn_bits = io_connPE_51_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_51_io_addressOut_ready = networkUnits_51_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_52_clock = clock;
  assign queues_52_reset = reset;
  assign queues_52_io_addressIn_valid = io_connPE_52_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_52_io_addressIn_bits = io_connPE_52_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_52_io_addressOut_ready = networkUnits_52_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_53_clock = clock;
  assign queues_53_reset = reset;
  assign queues_53_io_addressIn_valid = io_connPE_53_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_53_io_addressIn_bits = io_connPE_53_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_53_io_addressOut_ready = networkUnits_53_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_54_clock = clock;
  assign queues_54_reset = reset;
  assign queues_54_io_addressIn_valid = io_connPE_54_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_54_io_addressIn_bits = io_connPE_54_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_54_io_addressOut_ready = networkUnits_54_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_55_clock = clock;
  assign queues_55_reset = reset;
  assign queues_55_io_addressIn_valid = io_connPE_55_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_55_io_addressIn_bits = io_connPE_55_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_55_io_addressOut_ready = networkUnits_55_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_56_clock = clock;
  assign queues_56_reset = reset;
  assign queues_56_io_addressIn_valid = io_connPE_56_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_56_io_addressIn_bits = io_connPE_56_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_56_io_addressOut_ready = networkUnits_56_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_57_clock = clock;
  assign queues_57_reset = reset;
  assign queues_57_io_addressIn_valid = io_connPE_57_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_57_io_addressIn_bits = io_connPE_57_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_57_io_addressOut_ready = networkUnits_57_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_58_clock = clock;
  assign queues_58_reset = reset;
  assign queues_58_io_addressIn_valid = io_connPE_58_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_58_io_addressIn_bits = io_connPE_58_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_58_io_addressOut_ready = networkUnits_58_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_59_clock = clock;
  assign queues_59_reset = reset;
  assign queues_59_io_addressIn_valid = io_connPE_59_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_59_io_addressIn_bits = io_connPE_59_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_59_io_addressOut_ready = networkUnits_59_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_60_clock = clock;
  assign queues_60_reset = reset;
  assign queues_60_io_addressIn_valid = io_connPE_60_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_60_io_addressIn_bits = io_connPE_60_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_60_io_addressOut_ready = networkUnits_60_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_61_clock = clock;
  assign queues_61_reset = reset;
  assign queues_61_io_addressIn_valid = io_connPE_61_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_61_io_addressIn_bits = io_connPE_61_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_61_io_addressOut_ready = networkUnits_61_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_62_clock = clock;
  assign queues_62_reset = reset;
  assign queues_62_io_addressIn_valid = io_connPE_62_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_62_io_addressIn_bits = io_connPE_62_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_62_io_addressOut_ready = networkUnits_62_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
  assign queues_63_clock = clock;
  assign queues_63_reset = reset;
  assign queues_63_io_addressIn_valid = io_connPE_63_valid; // @[argRouteNetwork.scala 83:21]
  assign queues_63_io_addressIn_bits = io_connPE_63_bits; // @[argRouteNetwork.scala 83:21]
  assign queues_63_io_addressOut_ready = networkUnits_63_io_peAddress_ready; // @[argRouteNetwork.scala 92:38]
endmodule
module Queue_135(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram [0:15]; // @[Decoupled.scala 275:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 275:95]
  wire [3:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 275:95]
  wire [63:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 275:95]
  wire [63:0] ram_MPORT_data; // @[Decoupled.scala 275:95]
  wire [3:0] ram_MPORT_addr; // @[Decoupled.scala 275:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 275:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 275:95]
  reg [3:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [3:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 278:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 279:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 280:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 281:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 52:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 52:35]
  wire [3:0] _value_T_1 = enq_ptr_value + 4'h1; // @[Counter.scala 77:24]
  wire [3:0] _value_T_3 = deq_ptr_value + 4'h1; // @[Counter.scala 77:24]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 275:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 305:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 304:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 312:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 275:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 4'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 288:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 4'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 292:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 278:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 278:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 295:27]
      maybe_full <= do_enq; // @[Decoupled.scala 296:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_136(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram [0:15]; // @[Decoupled.scala 275:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 275:95]
  wire [3:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 275:95]
  wire [63:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 275:95]
  wire [63:0] ram_MPORT_data; // @[Decoupled.scala 275:95]
  wire [3:0] ram_MPORT_addr; // @[Decoupled.scala 275:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 275:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 275:95]
  reg [3:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [3:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 278:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 279:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 280:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 281:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 52:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 52:35]
  wire [3:0] _value_T_1 = enq_ptr_value + 4'h1; // @[Counter.scala 77:24]
  wire [3:0] _value_T_3 = deq_ptr_value + 4'h1; // @[Counter.scala 77:24]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 275:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 305:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 304:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 312:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 275:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 4'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 288:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 4'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 292:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 278:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 278:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 295:27]
      maybe_full <= do_enq; // @[Decoupled.scala 296:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module argRouteVirtServerV2(
  input          clock,
  input          reset,
  output         io_connNetwork_ready,
  input          io_connNetwork_valid,
  input  [63:0]  io_connNetwork_bits,
  input          io_connStealNtw_ctrl_serveStealReq_ready,
  output         io_connStealNtw_ctrl_serveStealReq_valid,
  input          io_connStealNtw_data_qOutTask_ready,
  output         io_connStealNtw_data_qOutTask_valid,
  output [255:0] io_connStealNtw_data_qOutTask_bits,
  input          io_read_address_ready,
  output         io_read_address_valid,
  output [63:0]  io_read_address_bits,
  output         io_read_data_ready,
  input          io_read_data_valid,
  input  [31:0]  io_read_data_bits,
  input          io_write_address_ready,
  output         io_write_address_valid,
  output [63:0]  io_write_address_bits,
  input          io_write_data_ready,
  output         io_write_data_valid,
  output [31:0]  io_write_data_bits,
  input          io_read_address_task_ready,
  output         io_read_address_task_valid,
  output [63:0]  io_read_address_task_bits,
  output         io_read_data_task_ready,
  input          io_read_data_task_valid,
  input  [31:0]  io_read_data_task_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [255:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  wire  addrNtwInQueue_clock; // @[argRouteServerV2.scala 48:32]
  wire  addrNtwInQueue_reset; // @[argRouteServerV2.scala 48:32]
  wire  addrNtwInQueue_io_enq_ready; // @[argRouteServerV2.scala 48:32]
  wire  addrNtwInQueue_io_enq_valid; // @[argRouteServerV2.scala 48:32]
  wire [63:0] addrNtwInQueue_io_enq_bits; // @[argRouteServerV2.scala 48:32]
  wire  addrNtwInQueue_io_deq_ready; // @[argRouteServerV2.scala 48:32]
  wire  addrNtwInQueue_io_deq_valid; // @[argRouteServerV2.scala 48:32]
  wire [63:0] addrNtwInQueue_io_deq_bits; // @[argRouteServerV2.scala 48:32]
  wire  addressesOfReadyTasks_clock; // @[argRouteServerV2.scala 53:39]
  wire  addressesOfReadyTasks_reset; // @[argRouteServerV2.scala 53:39]
  wire  addressesOfReadyTasks_io_enq_ready; // @[argRouteServerV2.scala 53:39]
  wire  addressesOfReadyTasks_io_enq_valid; // @[argRouteServerV2.scala 53:39]
  wire [63:0] addressesOfReadyTasks_io_enq_bits; // @[argRouteServerV2.scala 53:39]
  wire  addressesOfReadyTasks_io_deq_ready; // @[argRouteServerV2.scala 53:39]
  wire  addressesOfReadyTasks_io_deq_valid; // @[argRouteServerV2.scala 53:39]
  wire [63:0] addressesOfReadyTasks_io_deq_bits; // @[argRouteServerV2.scala 53:39]
  wire  readyTasksQueue_clock; // @[argRouteServerV2.scala 54:33]
  wire  readyTasksQueue_reset; // @[argRouteServerV2.scala 54:33]
  wire  readyTasksQueue_io_enq_ready; // @[argRouteServerV2.scala 54:33]
  wire  readyTasksQueue_io_enq_valid; // @[argRouteServerV2.scala 54:33]
  wire [255:0] readyTasksQueue_io_enq_bits; // @[argRouteServerV2.scala 54:33]
  wire  readyTasksQueue_io_deq_ready; // @[argRouteServerV2.scala 54:33]
  wire  readyTasksQueue_io_deq_valid; // @[argRouteServerV2.scala 54:33]
  wire [255:0] readyTasksQueue_io_deq_bits; // @[argRouteServerV2.scala 54:33]
  wire [4:0] readyTasksQueue_io_count; // @[argRouteServerV2.scala 54:33]
  reg [3:0] counterStateReg; // @[argRouteServerV2.scala 78:46]
  reg [63:0] counterReg; // @[argRouteServerV2.scala 79:46]
  reg [63:0] currReadAddr; // @[argRouteServerV2.scala 80:46]
  reg [63:0] counterAddr; // @[argRouteServerV2.scala 81:46]
  reg [63:0] addrMask; // @[argRouteServerV2.scala 82:46]
  wire  _T = counterStateReg == 4'h1; // @[argRouteServerV2.scala 103:26]
  wire [63:0] _counterAddr_T = addrNtwInQueue_io_deq_bits & addrMask; // @[argRouteServerV2.scala 106:55]
  wire  _T_1 = counterStateReg == 4'h2; // @[argRouteServerV2.scala 108:32]
  wire  _T_2 = counterStateReg == 4'h3; // @[argRouteServerV2.scala 112:32]
  wire [63:0] _currReadAddr_T_1 = counterAddr + 64'h4; // @[argRouteServerV2.scala 116:41]
  wire [31:0] _counterReg_T_1 = io_read_data_bits - 32'h1; // @[argRouteServerV2.scala 119:45]
  wire [63:0] _GEN_3 = io_read_data_valid ? {{32'd0}, _counterReg_T_1} : counterReg; // @[argRouteServerV2.scala 118:39 119:24 79:46]
  wire [3:0] _GEN_4 = io_read_data_valid ? 4'h4 : counterStateReg; // @[argRouteServerV2.scala 118:39 120:29 78:46]
  wire [63:0] _GEN_5 = io_read_data_valid & io_read_data_bits == 32'h1 ? _currReadAddr_T_1 : currReadAddr; // @[argRouteServerV2.scala 113:62 116:26 80:46]
  wire [3:0] _GEN_6 = io_read_data_valid & io_read_data_bits == 32'h1 ? 4'h7 : _GEN_4; // @[argRouteServerV2.scala 113:62 117:29]
  wire [63:0] _GEN_7 = io_read_data_valid & io_read_data_bits == 32'h1 ? counterReg : _GEN_3; // @[argRouteServerV2.scala 113:62 79:46]
  wire  _T_5 = counterStateReg == 4'h4; // @[argRouteServerV2.scala 122:32]
  wire [3:0] _GEN_8 = io_write_address_ready ? 4'h5 : counterStateReg; // @[argRouteServerV2.scala 123:37 124:29 78:46]
  wire  _T_6 = counterStateReg == 4'h5; // @[argRouteServerV2.scala 126:32]
  wire [3:0] _GEN_9 = io_write_data_ready ? 4'h1 : counterStateReg; // @[argRouteServerV2.scala 127:34 128:29 78:46]
  wire  _T_7 = counterStateReg == 4'h7; // @[argRouteServerV2.scala 130:32]
  wire [3:0] _GEN_10 = addressesOfReadyTasks_io_enq_ready ? 4'h1 : counterStateReg; // @[argRouteServerV2.scala 131:49 132:29 78:46]
  wire [3:0] _GEN_11 = counterStateReg == 4'h7 ? _GEN_10 : counterStateReg; // @[argRouteServerV2.scala 130:58 78:46]
  wire [3:0] _GEN_12 = counterStateReg == 4'h5 ? _GEN_9 : _GEN_11; // @[argRouteServerV2.scala 126:60]
  wire [3:0] _GEN_13 = counterStateReg == 4'h4 ? _GEN_8 : _GEN_12; // @[argRouteServerV2.scala 122:60]
  wire  _GEN_26 = _T_6 ? 1'h0 : _T_7; // @[argRouteServerV2.scala 144:60 88:40]
  wire  _GEN_28 = _T_5 ? 1'h0 : _T_6; // @[argRouteServerV2.scala 142:60 97:27]
  wire  _GEN_29 = _T_5 ? 1'h0 : _GEN_26; // @[argRouteServerV2.scala 142:60 88:40]
  wire  _GEN_31 = _T_2 ? 1'h0 : _T_5; // @[argRouteServerV2.scala 140:59 96:27]
  wire  _GEN_32 = _T_2 ? 1'h0 : _GEN_28; // @[argRouteServerV2.scala 140:59 97:27]
  wire  _GEN_33 = _T_2 ? 1'h0 : _GEN_29; // @[argRouteServerV2.scala 140:59 88:40]
  wire  _GEN_35 = _T_1 ? 1'h0 : _T_2; // @[argRouteServerV2.scala 138:59 98:27]
  wire  _GEN_36 = _T_1 ? 1'h0 : _GEN_31; // @[argRouteServerV2.scala 138:59 96:27]
  wire  _GEN_37 = _T_1 ? 1'h0 : _GEN_32; // @[argRouteServerV2.scala 138:59 97:27]
  wire  _GEN_38 = _T_1 ? 1'h0 : _GEN_33; // @[argRouteServerV2.scala 138:59 88:40]
  reg [3:0] taskReadAddressStateReg; // @[argRouteServerV2.scala 159:50]
  reg [63:0] taskAddr; // @[argRouteServerV2.scala 160:50]
  wire  _T_14 = taskReadAddressStateReg == 4'h6; // @[argRouteServerV2.scala 170:34]
  wire  _T_15 = taskReadAddressStateReg == 4'h8; // @[argRouteServerV2.scala 176:40]
  wire [63:0] _GEN_52 = _T_15 ? taskAddr : 64'h0; // @[argRouteServerV2.scala 167:32 193:71 195:36]
  reg [3:0] taskReadStateReg; // @[argRouteServerV2.scala 206:43]
  reg [2:0] taskReadCount; // @[argRouteServerV2.scala 207:43]
  reg [31:0] taskRegisters_0; // @[argRouteServerV2.scala 208:40]
  reg [31:0] taskRegisters_1; // @[argRouteServerV2.scala 208:40]
  reg [31:0] taskRegisters_2; // @[argRouteServerV2.scala 208:40]
  reg [31:0] taskRegisters_3; // @[argRouteServerV2.scala 208:40]
  reg [31:0] taskRegisters_4; // @[argRouteServerV2.scala 208:40]
  reg [31:0] taskRegisters_5; // @[argRouteServerV2.scala 208:40]
  reg [31:0] taskRegisters_6; // @[argRouteServerV2.scala 208:40]
  reg [31:0] taskRegisters_7; // @[argRouteServerV2.scala 208:40]
  wire [223:0] _readyTasksQueue_io_enq_bits_T_5 = {taskRegisters_0,taskRegisters_1,taskRegisters_2,taskRegisters_3,
    taskRegisters_4,taskRegisters_5,taskRegisters_6}; // @[Cat.scala 33:92]
  wire  _T_18 = taskReadStateReg == 4'h9; // @[argRouteServerV2.scala 217:27]
  wire [2:0] _T_20 = taskReadCount - 3'h1; // @[argRouteServerV2.scala 220:40]
  wire  _T_25 = taskReadStateReg == 4'ha; // @[argRouteServerV2.scala 228:33]
  reg [31:0] tasksGivenAwayCount; // @[argRouteServerV2.scala 247:48]
  reg [255:0] taskReg; // @[argRouteServerV2.scala 248:34]
  reg [3:0] taskWriteStateReg; // @[argRouteServerV2.scala 249:44]
  wire  _T_28 = taskWriteStateReg == 4'hb; // @[argRouteServerV2.scala 258:28]
  wire  _T_29 = taskWriteStateReg == 4'hc; // @[argRouteServerV2.scala 263:34]
  wire [31:0] _tasksGivenAwayCount_T_1 = tasksGivenAwayCount + 32'h1; // @[argRouteServerV2.scala 266:56]
  wire [31:0] _GEN_94 = io_connStealNtw_data_qOutTask_ready ? _tasksGivenAwayCount_T_1 : tasksGivenAwayCount; // @[argRouteServerV2.scala 264:50 266:33 247:48]
  wire [31:0] _GEN_96 = taskWriteStateReg == 4'hc ? _GEN_94 : tasksGivenAwayCount; // @[argRouteServerV2.scala 247:48 263:57]
  wire [31:0] _GEN_99 = taskWriteStateReg == 4'hb ? tasksGivenAwayCount : _GEN_96; // @[argRouteServerV2.scala 247:48 258:57]
  wire [31:0] _tasksGivenAwayCount_T_3 = tasksGivenAwayCount - 32'h1; // @[argRouteServerV2.scala 293:56]
  wire [70:0] _GEN_106 = reset ? 71'h0 : 71'h1fffffffffffffffe0; // @[argRouteServerV2.scala 82:{46,46} 83:37]
  Queue_135 addrNtwInQueue ( // @[argRouteServerV2.scala 48:32]
    .clock(addrNtwInQueue_clock),
    .reset(addrNtwInQueue_reset),
    .io_enq_ready(addrNtwInQueue_io_enq_ready),
    .io_enq_valid(addrNtwInQueue_io_enq_valid),
    .io_enq_bits(addrNtwInQueue_io_enq_bits),
    .io_deq_ready(addrNtwInQueue_io_deq_ready),
    .io_deq_valid(addrNtwInQueue_io_deq_valid),
    .io_deq_bits(addrNtwInQueue_io_deq_bits)
  );
  Queue_136 addressesOfReadyTasks ( // @[argRouteServerV2.scala 53:39]
    .clock(addressesOfReadyTasks_clock),
    .reset(addressesOfReadyTasks_reset),
    .io_enq_ready(addressesOfReadyTasks_io_enq_ready),
    .io_enq_valid(addressesOfReadyTasks_io_enq_valid),
    .io_enq_bits(addressesOfReadyTasks_io_enq_bits),
    .io_deq_ready(addressesOfReadyTasks_io_deq_ready),
    .io_deq_valid(addressesOfReadyTasks_io_deq_valid),
    .io_deq_bits(addressesOfReadyTasks_io_deq_bits)
  );
  Queue_3 readyTasksQueue ( // @[argRouteServerV2.scala 54:33]
    .clock(readyTasksQueue_clock),
    .reset(readyTasksQueue_reset),
    .io_enq_ready(readyTasksQueue_io_enq_ready),
    .io_enq_valid(readyTasksQueue_io_enq_valid),
    .io_enq_bits(readyTasksQueue_io_enq_bits),
    .io_deq_ready(readyTasksQueue_io_deq_ready),
    .io_deq_valid(readyTasksQueue_io_deq_valid),
    .io_deq_bits(readyTasksQueue_io_deq_bits),
    .io_count(readyTasksQueue_io_count)
  );
  assign io_connNetwork_ready = addrNtwInQueue_io_enq_ready; // @[argRouteServerV2.scala 57:27]
  assign io_connStealNtw_ctrl_serveStealReq_valid = tasksGivenAwayCount > 32'h0 & taskWriteStateReg != 4'hc; // @[argRouteServerV2.scala 290:36]
  assign io_connStealNtw_data_qOutTask_valid = _T_28 ? 1'h0 : _T_29; // @[argRouteServerV2.scala 256:46 270:57]
  assign io_connStealNtw_data_qOutTask_bits = taskReg; // @[argRouteServerV2.scala 254:46]
  assign io_read_address_valid = _T ? 1'h0 : _T_1; // @[argRouteServerV2.scala 136:48 95:27]
  assign io_read_address_bits = counterAddr; // @[argRouteServerV2.scala 92:27]
  assign io_read_data_ready = _T ? 1'h0 : _GEN_35; // @[argRouteServerV2.scala 136:48 98:27]
  assign io_write_address_valid = _T ? 1'h0 : _GEN_36; // @[argRouteServerV2.scala 136:48 96:27]
  assign io_write_address_bits = counterAddr; // @[argRouteServerV2.scala 93:27]
  assign io_write_data_valid = _T ? 1'h0 : _GEN_37; // @[argRouteServerV2.scala 136:48 97:27]
  assign io_write_data_bits = counterReg[31:0]; // @[argRouteServerV2.scala 94:27]
  assign io_read_address_task_valid = _T_14 ? 1'h0 : _T_15; // @[argRouteServerV2.scala 168:32 191:60]
  assign io_read_address_task_bits = _T_14 ? 64'h0 : _GEN_52; // @[argRouteServerV2.scala 167:32 191:60]
  assign io_read_data_task_ready = taskReadStateReg == 4'h9; // @[argRouteServerV2.scala 235:27]
  assign addrNtwInQueue_clock = clock;
  assign addrNtwInQueue_reset = reset;
  assign addrNtwInQueue_io_enq_valid = io_connNetwork_valid; // @[argRouteServerV2.scala 57:27]
  assign addrNtwInQueue_io_enq_bits = io_connNetwork_bits; // @[argRouteServerV2.scala 57:27]
  assign addrNtwInQueue_io_deq_ready = counterStateReg == 4'h1; // @[argRouteServerV2.scala 136:26]
  assign addressesOfReadyTasks_clock = clock;
  assign addressesOfReadyTasks_reset = reset;
  assign addressesOfReadyTasks_io_enq_valid = _T ? 1'h0 : _GEN_38; // @[argRouteServerV2.scala 136:48 88:40]
  assign addressesOfReadyTasks_io_enq_bits = currReadAddr; // @[argRouteServerV2.scala 89:40]
  assign addressesOfReadyTasks_io_deq_ready = taskReadAddressStateReg == 4'h6; // @[argRouteServerV2.scala 191:34]
  assign readyTasksQueue_clock = clock;
  assign readyTasksQueue_reset = reset;
  assign readyTasksQueue_io_enq_valid = _T_18 ? 1'h0 : _T_25; // @[argRouteServerV2.scala 211:34 235:46]
  assign readyTasksQueue_io_enq_bits = {_readyTasksQueue_io_enq_bits_T_5,taskRegisters_7}; // @[Cat.scala 33:92]
  assign readyTasksQueue_io_deq_ready = taskWriteStateReg == 4'hb; // @[argRouteServerV2.scala 270:28]
  always @(posedge clock) begin
    if (reset) begin // @[argRouteServerV2.scala 78:46]
      counterStateReg <= 4'h1; // @[argRouteServerV2.scala 78:46]
    end else if (counterStateReg == 4'h1) begin // @[argRouteServerV2.scala 103:48]
      if (addrNtwInQueue_io_deq_valid) begin // @[argRouteServerV2.scala 104:42]
        counterStateReg <= 4'h2; // @[argRouteServerV2.scala 105:32]
      end
    end else if (counterStateReg == 4'h2) begin // @[argRouteServerV2.scala 108:59]
      if (io_read_address_ready) begin // @[argRouteServerV2.scala 109:36]
        counterStateReg <= 4'h3; // @[argRouteServerV2.scala 110:29]
      end
    end else if (counterStateReg == 4'h3) begin // @[argRouteServerV2.scala 112:59]
      counterStateReg <= _GEN_6;
    end else begin
      counterStateReg <= _GEN_13;
    end
    if (reset) begin // @[argRouteServerV2.scala 79:46]
      counterReg <= 64'h0; // @[argRouteServerV2.scala 79:46]
    end else if (!(counterStateReg == 4'h1)) begin // @[argRouteServerV2.scala 103:48]
      if (!(counterStateReg == 4'h2)) begin // @[argRouteServerV2.scala 108:59]
        if (counterStateReg == 4'h3) begin // @[argRouteServerV2.scala 112:59]
          counterReg <= _GEN_7;
        end
      end
    end
    if (reset) begin // @[argRouteServerV2.scala 80:46]
      currReadAddr <= 64'h0; // @[argRouteServerV2.scala 80:46]
    end else if (!(counterStateReg == 4'h1)) begin // @[argRouteServerV2.scala 103:48]
      if (!(counterStateReg == 4'h2)) begin // @[argRouteServerV2.scala 108:59]
        if (counterStateReg == 4'h3) begin // @[argRouteServerV2.scala 112:59]
          currReadAddr <= _GEN_5;
        end
      end
    end
    if (reset) begin // @[argRouteServerV2.scala 81:46]
      counterAddr <= 64'h0; // @[argRouteServerV2.scala 81:46]
    end else if (counterStateReg == 4'h1) begin // @[argRouteServerV2.scala 103:48]
      if (addrNtwInQueue_io_deq_valid) begin // @[argRouteServerV2.scala 104:42]
        counterAddr <= _counterAddr_T; // @[argRouteServerV2.scala 106:25]
      end
    end
    addrMask <= _GEN_106[63:0]; // @[argRouteServerV2.scala 82:{46,46} 83:37]
    if (reset) begin // @[argRouteServerV2.scala 159:50]
      taskReadAddressStateReg <= 4'h6; // @[argRouteServerV2.scala 159:50]
    end else if (taskReadAddressStateReg == 4'h6) begin // @[argRouteServerV2.scala 170:60]
      if (addressesOfReadyTasks_io_deq_valid) begin // @[argRouteServerV2.scala 171:49]
        taskReadAddressStateReg <= 4'h8; // @[argRouteServerV2.scala 172:37]
      end
    end else if (taskReadAddressStateReg == 4'h8) begin // @[argRouteServerV2.scala 176:71]
      if (io_read_address_task_ready) begin // @[argRouteServerV2.scala 186:41]
        taskReadAddressStateReg <= 4'h6; // @[argRouteServerV2.scala 187:45]
      end
    end
    if (reset) begin // @[argRouteServerV2.scala 160:50]
      taskAddr <= 64'h0; // @[argRouteServerV2.scala 160:50]
    end else if (taskReadAddressStateReg == 4'h6) begin // @[argRouteServerV2.scala 170:60]
      if (addressesOfReadyTasks_io_deq_valid) begin // @[argRouteServerV2.scala 171:49]
        taskAddr <= addressesOfReadyTasks_io_deq_bits; // @[argRouteServerV2.scala 173:22]
      end
    end
    if (reset) begin // @[argRouteServerV2.scala 206:43]
      taskReadStateReg <= 4'h9; // @[argRouteServerV2.scala 206:43]
    end else if (taskReadStateReg == 4'h9) begin // @[argRouteServerV2.scala 217:46]
      if (taskReadCount == 3'h1 & io_read_data_task_valid) begin // @[argRouteServerV2.scala 224:63]
        taskReadStateReg <= 4'ha; // @[argRouteServerV2.scala 225:38]
      end
    end else if (taskReadStateReg == 4'ha) begin // @[argRouteServerV2.scala 228:61]
      if (readyTasksQueue_io_enq_ready) begin // @[argRouteServerV2.scala 229:43]
        taskReadStateReg <= 4'h9; // @[argRouteServerV2.scala 230:30]
      end
    end
    if (reset) begin // @[argRouteServerV2.scala 207:43]
      taskReadCount <= 3'h7; // @[argRouteServerV2.scala 207:43]
    end else if (taskReadStateReg == 4'h9) begin // @[argRouteServerV2.scala 217:46]
      if (io_read_data_task_valid) begin // @[argRouteServerV2.scala 219:38]
        taskReadCount <= _T_20; // @[argRouteServerV2.scala 221:27]
      end
    end else if (taskReadStateReg == 4'ha) begin // @[argRouteServerV2.scala 228:61]
      if (readyTasksQueue_io_enq_ready) begin // @[argRouteServerV2.scala 229:43]
        taskReadCount <= 3'h7; // @[argRouteServerV2.scala 231:30]
      end
    end
    if (reset) begin // @[argRouteServerV2.scala 208:40]
      taskRegisters_0 <= 32'h0; // @[argRouteServerV2.scala 208:40]
    end else if (taskReadStateReg == 4'h9) begin // @[argRouteServerV2.scala 217:46]
      if (io_read_data_task_valid) begin // @[argRouteServerV2.scala 219:38]
        if (3'h0 == _T_20) begin // @[argRouteServerV2.scala 220:46]
          taskRegisters_0 <= io_read_data_task_bits; // @[argRouteServerV2.scala 220:46]
        end
      end
    end
    if (reset) begin // @[argRouteServerV2.scala 208:40]
      taskRegisters_1 <= 32'h0; // @[argRouteServerV2.scala 208:40]
    end else if (taskReadStateReg == 4'h9) begin // @[argRouteServerV2.scala 217:46]
      if (io_read_data_task_valid) begin // @[argRouteServerV2.scala 219:38]
        if (3'h1 == _T_20) begin // @[argRouteServerV2.scala 220:46]
          taskRegisters_1 <= io_read_data_task_bits; // @[argRouteServerV2.scala 220:46]
        end
      end
    end
    if (reset) begin // @[argRouteServerV2.scala 208:40]
      taskRegisters_2 <= 32'h0; // @[argRouteServerV2.scala 208:40]
    end else if (taskReadStateReg == 4'h9) begin // @[argRouteServerV2.scala 217:46]
      if (io_read_data_task_valid) begin // @[argRouteServerV2.scala 219:38]
        if (3'h2 == _T_20) begin // @[argRouteServerV2.scala 220:46]
          taskRegisters_2 <= io_read_data_task_bits; // @[argRouteServerV2.scala 220:46]
        end
      end
    end
    if (reset) begin // @[argRouteServerV2.scala 208:40]
      taskRegisters_3 <= 32'h0; // @[argRouteServerV2.scala 208:40]
    end else if (taskReadStateReg == 4'h9) begin // @[argRouteServerV2.scala 217:46]
      if (io_read_data_task_valid) begin // @[argRouteServerV2.scala 219:38]
        if (3'h3 == _T_20) begin // @[argRouteServerV2.scala 220:46]
          taskRegisters_3 <= io_read_data_task_bits; // @[argRouteServerV2.scala 220:46]
        end
      end
    end
    if (reset) begin // @[argRouteServerV2.scala 208:40]
      taskRegisters_4 <= 32'h0; // @[argRouteServerV2.scala 208:40]
    end else if (taskReadStateReg == 4'h9) begin // @[argRouteServerV2.scala 217:46]
      if (io_read_data_task_valid) begin // @[argRouteServerV2.scala 219:38]
        if (3'h4 == _T_20) begin // @[argRouteServerV2.scala 220:46]
          taskRegisters_4 <= io_read_data_task_bits; // @[argRouteServerV2.scala 220:46]
        end
      end
    end
    if (reset) begin // @[argRouteServerV2.scala 208:40]
      taskRegisters_5 <= 32'h0; // @[argRouteServerV2.scala 208:40]
    end else if (taskReadStateReg == 4'h9) begin // @[argRouteServerV2.scala 217:46]
      if (io_read_data_task_valid) begin // @[argRouteServerV2.scala 219:38]
        if (3'h5 == _T_20) begin // @[argRouteServerV2.scala 220:46]
          taskRegisters_5 <= io_read_data_task_bits; // @[argRouteServerV2.scala 220:46]
        end
      end
    end
    if (reset) begin // @[argRouteServerV2.scala 208:40]
      taskRegisters_6 <= 32'h0; // @[argRouteServerV2.scala 208:40]
    end else if (taskReadStateReg == 4'h9) begin // @[argRouteServerV2.scala 217:46]
      if (io_read_data_task_valid) begin // @[argRouteServerV2.scala 219:38]
        if (3'h6 == _T_20) begin // @[argRouteServerV2.scala 220:46]
          taskRegisters_6 <= io_read_data_task_bits; // @[argRouteServerV2.scala 220:46]
        end
      end
    end
    if (reset) begin // @[argRouteServerV2.scala 208:40]
      taskRegisters_7 <= 32'h0; // @[argRouteServerV2.scala 208:40]
    end else if (taskReadStateReg == 4'h9) begin // @[argRouteServerV2.scala 217:46]
      if (io_read_data_task_valid) begin // @[argRouteServerV2.scala 219:38]
        if (3'h7 == _T_20) begin // @[argRouteServerV2.scala 220:46]
          taskRegisters_7 <= io_read_data_task_bits; // @[argRouteServerV2.scala 220:46]
        end
      end
    end
    if (reset) begin // @[argRouteServerV2.scala 247:48]
      tasksGivenAwayCount <= 32'h0; // @[argRouteServerV2.scala 247:48]
    end else if (tasksGivenAwayCount > 32'h0 & taskWriteStateReg != 4'hc) begin // @[argRouteServerV2.scala 290:80]
      if (io_connStealNtw_ctrl_serveStealReq_ready) begin // @[argRouteServerV2.scala 292:55]
        tasksGivenAwayCount <= _tasksGivenAwayCount_T_3; // @[argRouteServerV2.scala 293:33]
      end else begin
        tasksGivenAwayCount <= _GEN_99;
      end
    end else begin
      tasksGivenAwayCount <= _GEN_99;
    end
    if (reset) begin // @[argRouteServerV2.scala 248:34]
      taskReg <= 256'h0; // @[argRouteServerV2.scala 248:34]
    end else if (taskWriteStateReg == 4'hb) begin // @[argRouteServerV2.scala 258:57]
      if (readyTasksQueue_io_deq_valid) begin // @[argRouteServerV2.scala 259:43]
        taskReg <= readyTasksQueue_io_deq_bits; // @[argRouteServerV2.scala 261:21]
      end
    end
    if (reset) begin // @[argRouteServerV2.scala 249:44]
      taskWriteStateReg <= 4'hb; // @[argRouteServerV2.scala 249:44]
    end else if (taskWriteStateReg == 4'hb) begin // @[argRouteServerV2.scala 258:57]
      if (readyTasksQueue_io_deq_valid) begin // @[argRouteServerV2.scala 259:43]
        taskWriteStateReg <= 4'hc; // @[argRouteServerV2.scala 260:31]
      end
    end else if (taskWriteStateReg == 4'hc) begin // @[argRouteServerV2.scala 263:57]
      if (io_connStealNtw_data_qOutTask_ready) begin // @[argRouteServerV2.scala 264:50]
        taskWriteStateReg <= 4'hb; // @[argRouteServerV2.scala 265:31]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counterStateReg = _RAND_0[3:0];
  _RAND_1 = {2{`RANDOM}};
  counterReg = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  currReadAddr = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  counterAddr = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  addrMask = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  taskReadAddressStateReg = _RAND_5[3:0];
  _RAND_6 = {2{`RANDOM}};
  taskAddr = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  taskReadStateReg = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  taskReadCount = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  taskRegisters_0 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  taskRegisters_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  taskRegisters_2 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  taskRegisters_3 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  taskRegisters_4 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  taskRegisters_5 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  taskRegisters_6 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  taskRegisters_7 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  tasksGivenAwayCount = _RAND_17[31:0];
  _RAND_18 = {8{`RANDOM}};
  taskReg = _RAND_18[255:0];
  _RAND_19 = {1{`RANDOM}};
  taskWriteStateReg = _RAND_19[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module readyValidMem_2(
  input         clock,
  input         reset,
  output        io_read_address_ready,
  input         io_read_address_valid,
  input  [63:0] io_read_address_bits,
  input         io_read_data_ready,
  output        io_read_data_valid,
  output [31:0] io_read_data_bits,
  output        io_write_address_ready,
  input         io_write_address_valid,
  input  [63:0] io_write_address_bits,
  output        io_write_data_ready,
  input         io_write_data_valid,
  input  [31:0] io_write_data_bits,
  input         axi_ARREADY,
  output        axi_ARVALID,
  output [63:0] axi_ARADDR,
  output        axi_RREADY,
  input         axi_RVALID,
  input  [31:0] axi_RDATA,
  input         axi_AWREADY,
  output        axi_AWVALID,
  output [63:0] axi_AWADDR,
  input         axi_WREADY,
  output        axi_WVALID,
  output [31:0] axi_WDATA,
  input         axi_BVALID
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] writeDataDone; // @[readyValidMem.scala 47:30]
  reg  writeHandshakeDetector; // @[readyValidMem.scala 49:39]
  wire  _T_2 = writeDataDone == 2'h1; // @[readyValidMem.scala 100:32]
  wire  _GEN_2 = axi_BVALID ? 1'h0 : writeHandshakeDetector; // @[readyValidMem.scala 107:34 108:34 49:39]
  wire  _GEN_4 = io_write_data_valid & axi_WREADY & ~writeHandshakeDetector | _GEN_2; // @[readyValidMem.scala 104:82 106:34]
  assign io_read_address_ready = axi_ARREADY; // @[readyValidMem.scala 155:31]
  assign io_read_data_valid = axi_RVALID; // @[readyValidMem.scala 171:31]
  assign io_read_data_bits = axi_RDATA; // @[readyValidMem.scala 172:31]
  assign io_write_address_ready = axi_AWREADY; // @[readyValidMem.scala 143:32]
  assign io_write_data_ready = _T_2 & axi_BVALID; // @[readyValidMem.scala 111:62]
  assign axi_ARVALID = io_read_address_valid; // @[readyValidMem.scala 153:31]
  assign axi_ARADDR = io_read_address_bits; // @[readyValidMem.scala 154:31]
  assign axi_RREADY = io_read_data_ready; // @[readyValidMem.scala 169:31]
  assign axi_AWVALID = io_write_address_valid; // @[readyValidMem.scala 116:28]
  assign axi_AWADDR = io_write_address_bits; // @[readyValidMem.scala 117:28]
  assign axi_WVALID = io_write_data_valid & axi_WREADY & ~writeHandshakeDetector; // @[readyValidMem.scala 104:55]
  assign axi_WDATA = io_write_data_bits; // @[readyValidMem.scala 130:28]
  always @(posedge clock) begin
    if (reset) begin // @[readyValidMem.scala 47:30]
      writeDataDone <= 2'h0; // @[readyValidMem.scala 47:30]
    end else if (writeDataDone == 2'h0 & axi_WREADY) begin // @[readyValidMem.scala 98:53]
      writeDataDone <= 2'h1; // @[readyValidMem.scala 99:23]
    end else if (writeDataDone == 2'h1 & axi_BVALID) begin // @[readyValidMem.scala 100:59]
      writeDataDone <= 2'h0; // @[readyValidMem.scala 101:23]
    end
    if (reset) begin // @[readyValidMem.scala 49:39]
      writeHandshakeDetector <= 1'h0; // @[readyValidMem.scala 49:39]
    end else begin
      writeHandshakeDetector <= _GEN_4;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeDataDone = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  writeHandshakeDetector = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module readyValidMem_4(
  output        io_read_address_ready,
  input         io_read_address_valid,
  input  [63:0] io_read_address_bits,
  input         io_read_data_ready,
  output        io_read_data_valid,
  output [31:0] io_read_data_bits,
  input         axi_ARREADY,
  output        axi_ARVALID,
  output [63:0] axi_ARADDR,
  output        axi_RREADY,
  input         axi_RVALID,
  input  [31:0] axi_RDATA
);
  assign io_read_address_ready = axi_ARREADY; // @[readyValidMem.scala 155:31]
  assign io_read_data_valid = axi_RVALID; // @[readyValidMem.scala 171:31]
  assign io_read_data_bits = axi_RDATA; // @[readyValidMem.scala 172:31]
  assign axi_ARVALID = io_read_address_valid; // @[readyValidMem.scala 153:31]
  assign axi_ARADDR = io_read_address_bits; // @[readyValidMem.scala 154:31]
  assign axi_RREADY = io_read_data_ready; // @[readyValidMem.scala 169:31]
endmodule
module syncSide(
  input          clock,
  input          reset,
  output         io_addrIn_0_TREADY,
  input          io_addrIn_0_TVALID,
  input  [63:0]  io_addrIn_0_TDATA,
  output         io_addrIn_1_TREADY,
  input          io_addrIn_1_TVALID,
  input  [63:0]  io_addrIn_1_TDATA,
  output         io_addrIn_2_TREADY,
  input          io_addrIn_2_TVALID,
  input  [63:0]  io_addrIn_2_TDATA,
  output         io_addrIn_3_TREADY,
  input          io_addrIn_3_TVALID,
  input  [63:0]  io_addrIn_3_TDATA,
  output         io_addrIn_4_TREADY,
  input          io_addrIn_4_TVALID,
  input  [63:0]  io_addrIn_4_TDATA,
  output         io_addrIn_5_TREADY,
  input          io_addrIn_5_TVALID,
  input  [63:0]  io_addrIn_5_TDATA,
  output         io_addrIn_6_TREADY,
  input          io_addrIn_6_TVALID,
  input  [63:0]  io_addrIn_6_TDATA,
  output         io_addrIn_7_TREADY,
  input          io_addrIn_7_TVALID,
  input  [63:0]  io_addrIn_7_TDATA,
  output         io_addrIn_8_TREADY,
  input          io_addrIn_8_TVALID,
  input  [63:0]  io_addrIn_8_TDATA,
  output         io_addrIn_9_TREADY,
  input          io_addrIn_9_TVALID,
  input  [63:0]  io_addrIn_9_TDATA,
  output         io_addrIn_10_TREADY,
  input          io_addrIn_10_TVALID,
  input  [63:0]  io_addrIn_10_TDATA,
  output         io_addrIn_11_TREADY,
  input          io_addrIn_11_TVALID,
  input  [63:0]  io_addrIn_11_TDATA,
  output         io_addrIn_12_TREADY,
  input          io_addrIn_12_TVALID,
  input  [63:0]  io_addrIn_12_TDATA,
  output         io_addrIn_13_TREADY,
  input          io_addrIn_13_TVALID,
  input  [63:0]  io_addrIn_13_TDATA,
  output         io_addrIn_14_TREADY,
  input          io_addrIn_14_TVALID,
  input  [63:0]  io_addrIn_14_TDATA,
  output         io_addrIn_15_TREADY,
  input          io_addrIn_15_TVALID,
  input  [63:0]  io_addrIn_15_TDATA,
  output         io_addrIn_16_TREADY,
  input          io_addrIn_16_TVALID,
  input  [63:0]  io_addrIn_16_TDATA,
  output         io_addrIn_17_TREADY,
  input          io_addrIn_17_TVALID,
  input  [63:0]  io_addrIn_17_TDATA,
  output         io_addrIn_18_TREADY,
  input          io_addrIn_18_TVALID,
  input  [63:0]  io_addrIn_18_TDATA,
  output         io_addrIn_19_TREADY,
  input          io_addrIn_19_TVALID,
  input  [63:0]  io_addrIn_19_TDATA,
  output         io_addrIn_20_TREADY,
  input          io_addrIn_20_TVALID,
  input  [63:0]  io_addrIn_20_TDATA,
  output         io_addrIn_21_TREADY,
  input          io_addrIn_21_TVALID,
  input  [63:0]  io_addrIn_21_TDATA,
  output         io_addrIn_22_TREADY,
  input          io_addrIn_22_TVALID,
  input  [63:0]  io_addrIn_22_TDATA,
  output         io_addrIn_23_TREADY,
  input          io_addrIn_23_TVALID,
  input  [63:0]  io_addrIn_23_TDATA,
  output         io_addrIn_24_TREADY,
  input          io_addrIn_24_TVALID,
  input  [63:0]  io_addrIn_24_TDATA,
  output         io_addrIn_25_TREADY,
  input          io_addrIn_25_TVALID,
  input  [63:0]  io_addrIn_25_TDATA,
  output         io_addrIn_26_TREADY,
  input          io_addrIn_26_TVALID,
  input  [63:0]  io_addrIn_26_TDATA,
  output         io_addrIn_27_TREADY,
  input          io_addrIn_27_TVALID,
  input  [63:0]  io_addrIn_27_TDATA,
  output         io_addrIn_28_TREADY,
  input          io_addrIn_28_TVALID,
  input  [63:0]  io_addrIn_28_TDATA,
  output         io_addrIn_29_TREADY,
  input          io_addrIn_29_TVALID,
  input  [63:0]  io_addrIn_29_TDATA,
  output         io_addrIn_30_TREADY,
  input          io_addrIn_30_TVALID,
  input  [63:0]  io_addrIn_30_TDATA,
  output         io_addrIn_31_TREADY,
  input          io_addrIn_31_TVALID,
  input  [63:0]  io_addrIn_31_TDATA,
  output         io_addrIn_32_TREADY,
  input          io_addrIn_32_TVALID,
  input  [63:0]  io_addrIn_32_TDATA,
  output         io_addrIn_33_TREADY,
  input          io_addrIn_33_TVALID,
  input  [63:0]  io_addrIn_33_TDATA,
  output         io_addrIn_34_TREADY,
  input          io_addrIn_34_TVALID,
  input  [63:0]  io_addrIn_34_TDATA,
  output         io_addrIn_35_TREADY,
  input          io_addrIn_35_TVALID,
  input  [63:0]  io_addrIn_35_TDATA,
  output         io_addrIn_36_TREADY,
  input          io_addrIn_36_TVALID,
  input  [63:0]  io_addrIn_36_TDATA,
  output         io_addrIn_37_TREADY,
  input          io_addrIn_37_TVALID,
  input  [63:0]  io_addrIn_37_TDATA,
  output         io_addrIn_38_TREADY,
  input          io_addrIn_38_TVALID,
  input  [63:0]  io_addrIn_38_TDATA,
  output         io_addrIn_39_TREADY,
  input          io_addrIn_39_TVALID,
  input  [63:0]  io_addrIn_39_TDATA,
  output         io_addrIn_40_TREADY,
  input          io_addrIn_40_TVALID,
  input  [63:0]  io_addrIn_40_TDATA,
  output         io_addrIn_41_TREADY,
  input          io_addrIn_41_TVALID,
  input  [63:0]  io_addrIn_41_TDATA,
  output         io_addrIn_42_TREADY,
  input          io_addrIn_42_TVALID,
  input  [63:0]  io_addrIn_42_TDATA,
  output         io_addrIn_43_TREADY,
  input          io_addrIn_43_TVALID,
  input  [63:0]  io_addrIn_43_TDATA,
  output         io_addrIn_44_TREADY,
  input          io_addrIn_44_TVALID,
  input  [63:0]  io_addrIn_44_TDATA,
  output         io_addrIn_45_TREADY,
  input          io_addrIn_45_TVALID,
  input  [63:0]  io_addrIn_45_TDATA,
  output         io_addrIn_46_TREADY,
  input          io_addrIn_46_TVALID,
  input  [63:0]  io_addrIn_46_TDATA,
  output         io_addrIn_47_TREADY,
  input          io_addrIn_47_TVALID,
  input  [63:0]  io_addrIn_47_TDATA,
  output         io_addrIn_48_TREADY,
  input          io_addrIn_48_TVALID,
  input  [63:0]  io_addrIn_48_TDATA,
  output         io_addrIn_49_TREADY,
  input          io_addrIn_49_TVALID,
  input  [63:0]  io_addrIn_49_TDATA,
  output         io_addrIn_50_TREADY,
  input          io_addrIn_50_TVALID,
  input  [63:0]  io_addrIn_50_TDATA,
  output         io_addrIn_51_TREADY,
  input          io_addrIn_51_TVALID,
  input  [63:0]  io_addrIn_51_TDATA,
  output         io_addrIn_52_TREADY,
  input          io_addrIn_52_TVALID,
  input  [63:0]  io_addrIn_52_TDATA,
  output         io_addrIn_53_TREADY,
  input          io_addrIn_53_TVALID,
  input  [63:0]  io_addrIn_53_TDATA,
  output         io_addrIn_54_TREADY,
  input          io_addrIn_54_TVALID,
  input  [63:0]  io_addrIn_54_TDATA,
  output         io_addrIn_55_TREADY,
  input          io_addrIn_55_TVALID,
  input  [63:0]  io_addrIn_55_TDATA,
  output         io_addrIn_56_TREADY,
  input          io_addrIn_56_TVALID,
  input  [63:0]  io_addrIn_56_TDATA,
  output         io_addrIn_57_TREADY,
  input          io_addrIn_57_TVALID,
  input  [63:0]  io_addrIn_57_TDATA,
  output         io_addrIn_58_TREADY,
  input          io_addrIn_58_TVALID,
  input  [63:0]  io_addrIn_58_TDATA,
  output         io_addrIn_59_TREADY,
  input          io_addrIn_59_TVALID,
  input  [63:0]  io_addrIn_59_TDATA,
  output         io_addrIn_60_TREADY,
  input          io_addrIn_60_TVALID,
  input  [63:0]  io_addrIn_60_TDATA,
  output         io_addrIn_61_TREADY,
  input          io_addrIn_61_TVALID,
  input  [63:0]  io_addrIn_61_TDATA,
  output         io_addrIn_62_TREADY,
  input          io_addrIn_62_TVALID,
  input  [63:0]  io_addrIn_62_TDATA,
  output         io_addrIn_63_TREADY,
  input          io_addrIn_63_TVALID,
  input  [63:0]  io_addrIn_63_TDATA,
  input          io_axi_full_argRoute_0_ARREADY,
  output         io_axi_full_argRoute_0_ARVALID,
  output [63:0]  io_axi_full_argRoute_0_ARADDR,
  output         io_axi_full_argRoute_0_RREADY,
  input          io_axi_full_argRoute_0_RVALID,
  input  [31:0]  io_axi_full_argRoute_0_RDATA,
  input          io_axi_full_argRoute_0_AWREADY,
  output         io_axi_full_argRoute_0_AWVALID,
  output [63:0]  io_axi_full_argRoute_0_AWADDR,
  input          io_axi_full_argRoute_0_WREADY,
  output         io_axi_full_argRoute_0_WVALID,
  output [31:0]  io_axi_full_argRoute_0_WDATA,
  input          io_axi_full_argRoute_0_BVALID,
  input          io_axi_full_argRoute_1_ARREADY,
  output         io_axi_full_argRoute_1_ARVALID,
  output [63:0]  io_axi_full_argRoute_1_ARADDR,
  output         io_axi_full_argRoute_1_RREADY,
  input          io_axi_full_argRoute_1_RVALID,
  input  [31:0]  io_axi_full_argRoute_1_RDATA,
  input          io_axi_full_argRoute_1_AWREADY,
  output         io_axi_full_argRoute_1_AWVALID,
  output [63:0]  io_axi_full_argRoute_1_AWADDR,
  input          io_axi_full_argRoute_1_WREADY,
  output         io_axi_full_argRoute_1_WVALID,
  output [31:0]  io_axi_full_argRoute_1_WDATA,
  input          io_axi_full_argRoute_1_BVALID,
  input          io_axi_full_argRoute_2_ARREADY,
  output         io_axi_full_argRoute_2_ARVALID,
  output [63:0]  io_axi_full_argRoute_2_ARADDR,
  output         io_axi_full_argRoute_2_RREADY,
  input          io_axi_full_argRoute_2_RVALID,
  input  [31:0]  io_axi_full_argRoute_2_RDATA,
  input          io_axi_full_argRoute_3_ARREADY,
  output         io_axi_full_argRoute_3_ARVALID,
  output [63:0]  io_axi_full_argRoute_3_ARADDR,
  output         io_axi_full_argRoute_3_RREADY,
  input          io_axi_full_argRoute_3_RVALID,
  input  [31:0]  io_axi_full_argRoute_3_RDATA,
  input          connStealNtw_0_ctrl_serveStealReq_ready,
  output         connStealNtw_0_ctrl_serveStealReq_valid,
  input          connStealNtw_0_data_qOutTask_ready,
  output         connStealNtw_0_data_qOutTask_valid,
  output [255:0] connStealNtw_0_data_qOutTask_bits,
  input          connStealNtw_1_ctrl_serveStealReq_ready,
  output         connStealNtw_1_ctrl_serveStealReq_valid,
  input          connStealNtw_1_data_qOutTask_ready,
  output         connStealNtw_1_data_qOutTask_valid,
  output [255:0] connStealNtw_1_data_qOutTask_bits
);
  wire  argSide_clock; // @[syncSide.scala 46:25]
  wire  argSide_reset; // @[syncSide.scala 46:25]
  wire  argSide_io_connVAS_0_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connVAS_0_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connVAS_0_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connVAS_1_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connVAS_1_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connVAS_1_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_0_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_0_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_0_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_1_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_1_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_1_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_2_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_2_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_2_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_3_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_3_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_3_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_4_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_4_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_4_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_5_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_5_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_5_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_6_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_6_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_6_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_7_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_7_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_7_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_8_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_8_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_8_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_9_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_9_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_9_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_10_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_10_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_10_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_11_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_11_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_11_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_12_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_12_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_12_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_13_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_13_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_13_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_14_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_14_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_14_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_15_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_15_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_15_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_16_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_16_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_16_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_17_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_17_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_17_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_18_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_18_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_18_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_19_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_19_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_19_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_20_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_20_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_20_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_21_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_21_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_21_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_22_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_22_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_22_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_23_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_23_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_23_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_24_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_24_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_24_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_25_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_25_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_25_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_26_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_26_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_26_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_27_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_27_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_27_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_28_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_28_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_28_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_29_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_29_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_29_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_30_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_30_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_30_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_31_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_31_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_31_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_32_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_32_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_32_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_33_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_33_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_33_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_34_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_34_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_34_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_35_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_35_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_35_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_36_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_36_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_36_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_37_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_37_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_37_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_38_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_38_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_38_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_39_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_39_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_39_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_40_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_40_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_40_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_41_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_41_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_41_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_42_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_42_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_42_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_43_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_43_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_43_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_44_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_44_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_44_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_45_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_45_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_45_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_46_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_46_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_46_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_47_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_47_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_47_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_48_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_48_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_48_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_49_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_49_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_49_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_50_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_50_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_50_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_51_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_51_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_51_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_52_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_52_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_52_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_53_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_53_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_53_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_54_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_54_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_54_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_55_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_55_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_55_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_56_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_56_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_56_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_57_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_57_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_57_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_58_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_58_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_58_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_59_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_59_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_59_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_60_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_60_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_60_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_61_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_61_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_61_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_62_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_62_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_62_bits; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_63_ready; // @[syncSide.scala 46:25]
  wire  argSide_io_connPE_63_valid; // @[syncSide.scala 46:25]
  wire [63:0] argSide_io_connPE_63_bits; // @[syncSide.scala 46:25]
  wire  argRouteServers_0_clock; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_reset; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_io_connNetwork_ready; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_io_connNetwork_valid; // @[syncSide.scala 55:15]
  wire [63:0] argRouteServers_0_io_connNetwork_bits; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_io_connStealNtw_ctrl_serveStealReq_ready; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_io_connStealNtw_ctrl_serveStealReq_valid; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_io_connStealNtw_data_qOutTask_ready; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_io_connStealNtw_data_qOutTask_valid; // @[syncSide.scala 55:15]
  wire [255:0] argRouteServers_0_io_connStealNtw_data_qOutTask_bits; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_io_read_address_ready; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_io_read_address_valid; // @[syncSide.scala 55:15]
  wire [63:0] argRouteServers_0_io_read_address_bits; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_io_read_data_ready; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_io_read_data_valid; // @[syncSide.scala 55:15]
  wire [31:0] argRouteServers_0_io_read_data_bits; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_io_write_address_ready; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_io_write_address_valid; // @[syncSide.scala 55:15]
  wire [63:0] argRouteServers_0_io_write_address_bits; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_io_write_data_ready; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_io_write_data_valid; // @[syncSide.scala 55:15]
  wire [31:0] argRouteServers_0_io_write_data_bits; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_io_read_address_task_ready; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_io_read_address_task_valid; // @[syncSide.scala 55:15]
  wire [63:0] argRouteServers_0_io_read_address_task_bits; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_io_read_data_task_ready; // @[syncSide.scala 55:15]
  wire  argRouteServers_0_io_read_data_task_valid; // @[syncSide.scala 55:15]
  wire [31:0] argRouteServers_0_io_read_data_task_bits; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_clock; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_reset; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_io_connNetwork_ready; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_io_connNetwork_valid; // @[syncSide.scala 55:15]
  wire [63:0] argRouteServers_1_io_connNetwork_bits; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_io_connStealNtw_ctrl_serveStealReq_ready; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_io_connStealNtw_ctrl_serveStealReq_valid; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_io_connStealNtw_data_qOutTask_ready; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_io_connStealNtw_data_qOutTask_valid; // @[syncSide.scala 55:15]
  wire [255:0] argRouteServers_1_io_connStealNtw_data_qOutTask_bits; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_io_read_address_ready; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_io_read_address_valid; // @[syncSide.scala 55:15]
  wire [63:0] argRouteServers_1_io_read_address_bits; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_io_read_data_ready; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_io_read_data_valid; // @[syncSide.scala 55:15]
  wire [31:0] argRouteServers_1_io_read_data_bits; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_io_write_address_ready; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_io_write_address_valid; // @[syncSide.scala 55:15]
  wire [63:0] argRouteServers_1_io_write_address_bits; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_io_write_data_ready; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_io_write_data_valid; // @[syncSide.scala 55:15]
  wire [31:0] argRouteServers_1_io_write_data_bits; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_io_read_address_task_ready; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_io_read_address_task_valid; // @[syncSide.scala 55:15]
  wire [63:0] argRouteServers_1_io_read_address_task_bits; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_io_read_data_task_ready; // @[syncSide.scala 55:15]
  wire  argRouteServers_1_io_read_data_task_valid; // @[syncSide.scala 55:15]
  wire [31:0] argRouteServers_1_io_read_data_task_bits; // @[syncSide.scala 55:15]
  wire  argRouteRvm_0_clock; // @[syncSide.scala 65:67]
  wire  argRouteRvm_0_reset; // @[syncSide.scala 65:67]
  wire  argRouteRvm_0_io_read_address_ready; // @[syncSide.scala 65:67]
  wire  argRouteRvm_0_io_read_address_valid; // @[syncSide.scala 65:67]
  wire [63:0] argRouteRvm_0_io_read_address_bits; // @[syncSide.scala 65:67]
  wire  argRouteRvm_0_io_read_data_ready; // @[syncSide.scala 65:67]
  wire  argRouteRvm_0_io_read_data_valid; // @[syncSide.scala 65:67]
  wire [31:0] argRouteRvm_0_io_read_data_bits; // @[syncSide.scala 65:67]
  wire  argRouteRvm_0_io_write_address_ready; // @[syncSide.scala 65:67]
  wire  argRouteRvm_0_io_write_address_valid; // @[syncSide.scala 65:67]
  wire [63:0] argRouteRvm_0_io_write_address_bits; // @[syncSide.scala 65:67]
  wire  argRouteRvm_0_io_write_data_ready; // @[syncSide.scala 65:67]
  wire  argRouteRvm_0_io_write_data_valid; // @[syncSide.scala 65:67]
  wire [31:0] argRouteRvm_0_io_write_data_bits; // @[syncSide.scala 65:67]
  wire  argRouteRvm_0_axi_ARREADY; // @[syncSide.scala 65:67]
  wire  argRouteRvm_0_axi_ARVALID; // @[syncSide.scala 65:67]
  wire [63:0] argRouteRvm_0_axi_ARADDR; // @[syncSide.scala 65:67]
  wire  argRouteRvm_0_axi_RREADY; // @[syncSide.scala 65:67]
  wire  argRouteRvm_0_axi_RVALID; // @[syncSide.scala 65:67]
  wire [31:0] argRouteRvm_0_axi_RDATA; // @[syncSide.scala 65:67]
  wire  argRouteRvm_0_axi_AWREADY; // @[syncSide.scala 65:67]
  wire  argRouteRvm_0_axi_AWVALID; // @[syncSide.scala 65:67]
  wire [63:0] argRouteRvm_0_axi_AWADDR; // @[syncSide.scala 65:67]
  wire  argRouteRvm_0_axi_WREADY; // @[syncSide.scala 65:67]
  wire  argRouteRvm_0_axi_WVALID; // @[syncSide.scala 65:67]
  wire [31:0] argRouteRvm_0_axi_WDATA; // @[syncSide.scala 65:67]
  wire  argRouteRvm_0_axi_BVALID; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_clock; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_reset; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_io_read_address_ready; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_io_read_address_valid; // @[syncSide.scala 65:67]
  wire [63:0] argRouteRvm_1_io_read_address_bits; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_io_read_data_ready; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_io_read_data_valid; // @[syncSide.scala 65:67]
  wire [31:0] argRouteRvm_1_io_read_data_bits; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_io_write_address_ready; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_io_write_address_valid; // @[syncSide.scala 65:67]
  wire [63:0] argRouteRvm_1_io_write_address_bits; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_io_write_data_ready; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_io_write_data_valid; // @[syncSide.scala 65:67]
  wire [31:0] argRouteRvm_1_io_write_data_bits; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_axi_ARREADY; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_axi_ARVALID; // @[syncSide.scala 65:67]
  wire [63:0] argRouteRvm_1_axi_ARADDR; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_axi_RREADY; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_axi_RVALID; // @[syncSide.scala 65:67]
  wire [31:0] argRouteRvm_1_axi_RDATA; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_axi_AWREADY; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_axi_AWVALID; // @[syncSide.scala 65:67]
  wire [63:0] argRouteRvm_1_axi_AWADDR; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_axi_WREADY; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_axi_WVALID; // @[syncSide.scala 65:67]
  wire [31:0] argRouteRvm_1_axi_WDATA; // @[syncSide.scala 65:67]
  wire  argRouteRvm_1_axi_BVALID; // @[syncSide.scala 65:67]
  wire  argRouteRvmReadOnly_0_io_read_address_ready; // @[syncSide.scala 66:69]
  wire  argRouteRvmReadOnly_0_io_read_address_valid; // @[syncSide.scala 66:69]
  wire [63:0] argRouteRvmReadOnly_0_io_read_address_bits; // @[syncSide.scala 66:69]
  wire  argRouteRvmReadOnly_0_io_read_data_ready; // @[syncSide.scala 66:69]
  wire  argRouteRvmReadOnly_0_io_read_data_valid; // @[syncSide.scala 66:69]
  wire [31:0] argRouteRvmReadOnly_0_io_read_data_bits; // @[syncSide.scala 66:69]
  wire  argRouteRvmReadOnly_0_axi_ARREADY; // @[syncSide.scala 66:69]
  wire  argRouteRvmReadOnly_0_axi_ARVALID; // @[syncSide.scala 66:69]
  wire [63:0] argRouteRvmReadOnly_0_axi_ARADDR; // @[syncSide.scala 66:69]
  wire  argRouteRvmReadOnly_0_axi_RREADY; // @[syncSide.scala 66:69]
  wire  argRouteRvmReadOnly_0_axi_RVALID; // @[syncSide.scala 66:69]
  wire [31:0] argRouteRvmReadOnly_0_axi_RDATA; // @[syncSide.scala 66:69]
  wire  argRouteRvmReadOnly_1_io_read_address_ready; // @[syncSide.scala 66:69]
  wire  argRouteRvmReadOnly_1_io_read_address_valid; // @[syncSide.scala 66:69]
  wire [63:0] argRouteRvmReadOnly_1_io_read_address_bits; // @[syncSide.scala 66:69]
  wire  argRouteRvmReadOnly_1_io_read_data_ready; // @[syncSide.scala 66:69]
  wire  argRouteRvmReadOnly_1_io_read_data_valid; // @[syncSide.scala 66:69]
  wire [31:0] argRouteRvmReadOnly_1_io_read_data_bits; // @[syncSide.scala 66:69]
  wire  argRouteRvmReadOnly_1_axi_ARREADY; // @[syncSide.scala 66:69]
  wire  argRouteRvmReadOnly_1_axi_ARVALID; // @[syncSide.scala 66:69]
  wire [63:0] argRouteRvmReadOnly_1_axi_ARADDR; // @[syncSide.scala 66:69]
  wire  argRouteRvmReadOnly_1_axi_RREADY; // @[syncSide.scala 66:69]
  wire  argRouteRvmReadOnly_1_axi_RVALID; // @[syncSide.scala 66:69]
  wire [31:0] argRouteRvmReadOnly_1_axi_RDATA; // @[syncSide.scala 66:69]
  argRouteNetwork argSide ( // @[syncSide.scala 46:25]
    .clock(argSide_clock),
    .reset(argSide_reset),
    .io_connVAS_0_ready(argSide_io_connVAS_0_ready),
    .io_connVAS_0_valid(argSide_io_connVAS_0_valid),
    .io_connVAS_0_bits(argSide_io_connVAS_0_bits),
    .io_connVAS_1_ready(argSide_io_connVAS_1_ready),
    .io_connVAS_1_valid(argSide_io_connVAS_1_valid),
    .io_connVAS_1_bits(argSide_io_connVAS_1_bits),
    .io_connPE_0_ready(argSide_io_connPE_0_ready),
    .io_connPE_0_valid(argSide_io_connPE_0_valid),
    .io_connPE_0_bits(argSide_io_connPE_0_bits),
    .io_connPE_1_ready(argSide_io_connPE_1_ready),
    .io_connPE_1_valid(argSide_io_connPE_1_valid),
    .io_connPE_1_bits(argSide_io_connPE_1_bits),
    .io_connPE_2_ready(argSide_io_connPE_2_ready),
    .io_connPE_2_valid(argSide_io_connPE_2_valid),
    .io_connPE_2_bits(argSide_io_connPE_2_bits),
    .io_connPE_3_ready(argSide_io_connPE_3_ready),
    .io_connPE_3_valid(argSide_io_connPE_3_valid),
    .io_connPE_3_bits(argSide_io_connPE_3_bits),
    .io_connPE_4_ready(argSide_io_connPE_4_ready),
    .io_connPE_4_valid(argSide_io_connPE_4_valid),
    .io_connPE_4_bits(argSide_io_connPE_4_bits),
    .io_connPE_5_ready(argSide_io_connPE_5_ready),
    .io_connPE_5_valid(argSide_io_connPE_5_valid),
    .io_connPE_5_bits(argSide_io_connPE_5_bits),
    .io_connPE_6_ready(argSide_io_connPE_6_ready),
    .io_connPE_6_valid(argSide_io_connPE_6_valid),
    .io_connPE_6_bits(argSide_io_connPE_6_bits),
    .io_connPE_7_ready(argSide_io_connPE_7_ready),
    .io_connPE_7_valid(argSide_io_connPE_7_valid),
    .io_connPE_7_bits(argSide_io_connPE_7_bits),
    .io_connPE_8_ready(argSide_io_connPE_8_ready),
    .io_connPE_8_valid(argSide_io_connPE_8_valid),
    .io_connPE_8_bits(argSide_io_connPE_8_bits),
    .io_connPE_9_ready(argSide_io_connPE_9_ready),
    .io_connPE_9_valid(argSide_io_connPE_9_valid),
    .io_connPE_9_bits(argSide_io_connPE_9_bits),
    .io_connPE_10_ready(argSide_io_connPE_10_ready),
    .io_connPE_10_valid(argSide_io_connPE_10_valid),
    .io_connPE_10_bits(argSide_io_connPE_10_bits),
    .io_connPE_11_ready(argSide_io_connPE_11_ready),
    .io_connPE_11_valid(argSide_io_connPE_11_valid),
    .io_connPE_11_bits(argSide_io_connPE_11_bits),
    .io_connPE_12_ready(argSide_io_connPE_12_ready),
    .io_connPE_12_valid(argSide_io_connPE_12_valid),
    .io_connPE_12_bits(argSide_io_connPE_12_bits),
    .io_connPE_13_ready(argSide_io_connPE_13_ready),
    .io_connPE_13_valid(argSide_io_connPE_13_valid),
    .io_connPE_13_bits(argSide_io_connPE_13_bits),
    .io_connPE_14_ready(argSide_io_connPE_14_ready),
    .io_connPE_14_valid(argSide_io_connPE_14_valid),
    .io_connPE_14_bits(argSide_io_connPE_14_bits),
    .io_connPE_15_ready(argSide_io_connPE_15_ready),
    .io_connPE_15_valid(argSide_io_connPE_15_valid),
    .io_connPE_15_bits(argSide_io_connPE_15_bits),
    .io_connPE_16_ready(argSide_io_connPE_16_ready),
    .io_connPE_16_valid(argSide_io_connPE_16_valid),
    .io_connPE_16_bits(argSide_io_connPE_16_bits),
    .io_connPE_17_ready(argSide_io_connPE_17_ready),
    .io_connPE_17_valid(argSide_io_connPE_17_valid),
    .io_connPE_17_bits(argSide_io_connPE_17_bits),
    .io_connPE_18_ready(argSide_io_connPE_18_ready),
    .io_connPE_18_valid(argSide_io_connPE_18_valid),
    .io_connPE_18_bits(argSide_io_connPE_18_bits),
    .io_connPE_19_ready(argSide_io_connPE_19_ready),
    .io_connPE_19_valid(argSide_io_connPE_19_valid),
    .io_connPE_19_bits(argSide_io_connPE_19_bits),
    .io_connPE_20_ready(argSide_io_connPE_20_ready),
    .io_connPE_20_valid(argSide_io_connPE_20_valid),
    .io_connPE_20_bits(argSide_io_connPE_20_bits),
    .io_connPE_21_ready(argSide_io_connPE_21_ready),
    .io_connPE_21_valid(argSide_io_connPE_21_valid),
    .io_connPE_21_bits(argSide_io_connPE_21_bits),
    .io_connPE_22_ready(argSide_io_connPE_22_ready),
    .io_connPE_22_valid(argSide_io_connPE_22_valid),
    .io_connPE_22_bits(argSide_io_connPE_22_bits),
    .io_connPE_23_ready(argSide_io_connPE_23_ready),
    .io_connPE_23_valid(argSide_io_connPE_23_valid),
    .io_connPE_23_bits(argSide_io_connPE_23_bits),
    .io_connPE_24_ready(argSide_io_connPE_24_ready),
    .io_connPE_24_valid(argSide_io_connPE_24_valid),
    .io_connPE_24_bits(argSide_io_connPE_24_bits),
    .io_connPE_25_ready(argSide_io_connPE_25_ready),
    .io_connPE_25_valid(argSide_io_connPE_25_valid),
    .io_connPE_25_bits(argSide_io_connPE_25_bits),
    .io_connPE_26_ready(argSide_io_connPE_26_ready),
    .io_connPE_26_valid(argSide_io_connPE_26_valid),
    .io_connPE_26_bits(argSide_io_connPE_26_bits),
    .io_connPE_27_ready(argSide_io_connPE_27_ready),
    .io_connPE_27_valid(argSide_io_connPE_27_valid),
    .io_connPE_27_bits(argSide_io_connPE_27_bits),
    .io_connPE_28_ready(argSide_io_connPE_28_ready),
    .io_connPE_28_valid(argSide_io_connPE_28_valid),
    .io_connPE_28_bits(argSide_io_connPE_28_bits),
    .io_connPE_29_ready(argSide_io_connPE_29_ready),
    .io_connPE_29_valid(argSide_io_connPE_29_valid),
    .io_connPE_29_bits(argSide_io_connPE_29_bits),
    .io_connPE_30_ready(argSide_io_connPE_30_ready),
    .io_connPE_30_valid(argSide_io_connPE_30_valid),
    .io_connPE_30_bits(argSide_io_connPE_30_bits),
    .io_connPE_31_ready(argSide_io_connPE_31_ready),
    .io_connPE_31_valid(argSide_io_connPE_31_valid),
    .io_connPE_31_bits(argSide_io_connPE_31_bits),
    .io_connPE_32_ready(argSide_io_connPE_32_ready),
    .io_connPE_32_valid(argSide_io_connPE_32_valid),
    .io_connPE_32_bits(argSide_io_connPE_32_bits),
    .io_connPE_33_ready(argSide_io_connPE_33_ready),
    .io_connPE_33_valid(argSide_io_connPE_33_valid),
    .io_connPE_33_bits(argSide_io_connPE_33_bits),
    .io_connPE_34_ready(argSide_io_connPE_34_ready),
    .io_connPE_34_valid(argSide_io_connPE_34_valid),
    .io_connPE_34_bits(argSide_io_connPE_34_bits),
    .io_connPE_35_ready(argSide_io_connPE_35_ready),
    .io_connPE_35_valid(argSide_io_connPE_35_valid),
    .io_connPE_35_bits(argSide_io_connPE_35_bits),
    .io_connPE_36_ready(argSide_io_connPE_36_ready),
    .io_connPE_36_valid(argSide_io_connPE_36_valid),
    .io_connPE_36_bits(argSide_io_connPE_36_bits),
    .io_connPE_37_ready(argSide_io_connPE_37_ready),
    .io_connPE_37_valid(argSide_io_connPE_37_valid),
    .io_connPE_37_bits(argSide_io_connPE_37_bits),
    .io_connPE_38_ready(argSide_io_connPE_38_ready),
    .io_connPE_38_valid(argSide_io_connPE_38_valid),
    .io_connPE_38_bits(argSide_io_connPE_38_bits),
    .io_connPE_39_ready(argSide_io_connPE_39_ready),
    .io_connPE_39_valid(argSide_io_connPE_39_valid),
    .io_connPE_39_bits(argSide_io_connPE_39_bits),
    .io_connPE_40_ready(argSide_io_connPE_40_ready),
    .io_connPE_40_valid(argSide_io_connPE_40_valid),
    .io_connPE_40_bits(argSide_io_connPE_40_bits),
    .io_connPE_41_ready(argSide_io_connPE_41_ready),
    .io_connPE_41_valid(argSide_io_connPE_41_valid),
    .io_connPE_41_bits(argSide_io_connPE_41_bits),
    .io_connPE_42_ready(argSide_io_connPE_42_ready),
    .io_connPE_42_valid(argSide_io_connPE_42_valid),
    .io_connPE_42_bits(argSide_io_connPE_42_bits),
    .io_connPE_43_ready(argSide_io_connPE_43_ready),
    .io_connPE_43_valid(argSide_io_connPE_43_valid),
    .io_connPE_43_bits(argSide_io_connPE_43_bits),
    .io_connPE_44_ready(argSide_io_connPE_44_ready),
    .io_connPE_44_valid(argSide_io_connPE_44_valid),
    .io_connPE_44_bits(argSide_io_connPE_44_bits),
    .io_connPE_45_ready(argSide_io_connPE_45_ready),
    .io_connPE_45_valid(argSide_io_connPE_45_valid),
    .io_connPE_45_bits(argSide_io_connPE_45_bits),
    .io_connPE_46_ready(argSide_io_connPE_46_ready),
    .io_connPE_46_valid(argSide_io_connPE_46_valid),
    .io_connPE_46_bits(argSide_io_connPE_46_bits),
    .io_connPE_47_ready(argSide_io_connPE_47_ready),
    .io_connPE_47_valid(argSide_io_connPE_47_valid),
    .io_connPE_47_bits(argSide_io_connPE_47_bits),
    .io_connPE_48_ready(argSide_io_connPE_48_ready),
    .io_connPE_48_valid(argSide_io_connPE_48_valid),
    .io_connPE_48_bits(argSide_io_connPE_48_bits),
    .io_connPE_49_ready(argSide_io_connPE_49_ready),
    .io_connPE_49_valid(argSide_io_connPE_49_valid),
    .io_connPE_49_bits(argSide_io_connPE_49_bits),
    .io_connPE_50_ready(argSide_io_connPE_50_ready),
    .io_connPE_50_valid(argSide_io_connPE_50_valid),
    .io_connPE_50_bits(argSide_io_connPE_50_bits),
    .io_connPE_51_ready(argSide_io_connPE_51_ready),
    .io_connPE_51_valid(argSide_io_connPE_51_valid),
    .io_connPE_51_bits(argSide_io_connPE_51_bits),
    .io_connPE_52_ready(argSide_io_connPE_52_ready),
    .io_connPE_52_valid(argSide_io_connPE_52_valid),
    .io_connPE_52_bits(argSide_io_connPE_52_bits),
    .io_connPE_53_ready(argSide_io_connPE_53_ready),
    .io_connPE_53_valid(argSide_io_connPE_53_valid),
    .io_connPE_53_bits(argSide_io_connPE_53_bits),
    .io_connPE_54_ready(argSide_io_connPE_54_ready),
    .io_connPE_54_valid(argSide_io_connPE_54_valid),
    .io_connPE_54_bits(argSide_io_connPE_54_bits),
    .io_connPE_55_ready(argSide_io_connPE_55_ready),
    .io_connPE_55_valid(argSide_io_connPE_55_valid),
    .io_connPE_55_bits(argSide_io_connPE_55_bits),
    .io_connPE_56_ready(argSide_io_connPE_56_ready),
    .io_connPE_56_valid(argSide_io_connPE_56_valid),
    .io_connPE_56_bits(argSide_io_connPE_56_bits),
    .io_connPE_57_ready(argSide_io_connPE_57_ready),
    .io_connPE_57_valid(argSide_io_connPE_57_valid),
    .io_connPE_57_bits(argSide_io_connPE_57_bits),
    .io_connPE_58_ready(argSide_io_connPE_58_ready),
    .io_connPE_58_valid(argSide_io_connPE_58_valid),
    .io_connPE_58_bits(argSide_io_connPE_58_bits),
    .io_connPE_59_ready(argSide_io_connPE_59_ready),
    .io_connPE_59_valid(argSide_io_connPE_59_valid),
    .io_connPE_59_bits(argSide_io_connPE_59_bits),
    .io_connPE_60_ready(argSide_io_connPE_60_ready),
    .io_connPE_60_valid(argSide_io_connPE_60_valid),
    .io_connPE_60_bits(argSide_io_connPE_60_bits),
    .io_connPE_61_ready(argSide_io_connPE_61_ready),
    .io_connPE_61_valid(argSide_io_connPE_61_valid),
    .io_connPE_61_bits(argSide_io_connPE_61_bits),
    .io_connPE_62_ready(argSide_io_connPE_62_ready),
    .io_connPE_62_valid(argSide_io_connPE_62_valid),
    .io_connPE_62_bits(argSide_io_connPE_62_bits),
    .io_connPE_63_ready(argSide_io_connPE_63_ready),
    .io_connPE_63_valid(argSide_io_connPE_63_valid),
    .io_connPE_63_bits(argSide_io_connPE_63_bits)
  );
  argRouteVirtServerV2 argRouteServers_0 ( // @[syncSide.scala 55:15]
    .clock(argRouteServers_0_clock),
    .reset(argRouteServers_0_reset),
    .io_connNetwork_ready(argRouteServers_0_io_connNetwork_ready),
    .io_connNetwork_valid(argRouteServers_0_io_connNetwork_valid),
    .io_connNetwork_bits(argRouteServers_0_io_connNetwork_bits),
    .io_connStealNtw_ctrl_serveStealReq_ready(argRouteServers_0_io_connStealNtw_ctrl_serveStealReq_ready),
    .io_connStealNtw_ctrl_serveStealReq_valid(argRouteServers_0_io_connStealNtw_ctrl_serveStealReq_valid),
    .io_connStealNtw_data_qOutTask_ready(argRouteServers_0_io_connStealNtw_data_qOutTask_ready),
    .io_connStealNtw_data_qOutTask_valid(argRouteServers_0_io_connStealNtw_data_qOutTask_valid),
    .io_connStealNtw_data_qOutTask_bits(argRouteServers_0_io_connStealNtw_data_qOutTask_bits),
    .io_read_address_ready(argRouteServers_0_io_read_address_ready),
    .io_read_address_valid(argRouteServers_0_io_read_address_valid),
    .io_read_address_bits(argRouteServers_0_io_read_address_bits),
    .io_read_data_ready(argRouteServers_0_io_read_data_ready),
    .io_read_data_valid(argRouteServers_0_io_read_data_valid),
    .io_read_data_bits(argRouteServers_0_io_read_data_bits),
    .io_write_address_ready(argRouteServers_0_io_write_address_ready),
    .io_write_address_valid(argRouteServers_0_io_write_address_valid),
    .io_write_address_bits(argRouteServers_0_io_write_address_bits),
    .io_write_data_ready(argRouteServers_0_io_write_data_ready),
    .io_write_data_valid(argRouteServers_0_io_write_data_valid),
    .io_write_data_bits(argRouteServers_0_io_write_data_bits),
    .io_read_address_task_ready(argRouteServers_0_io_read_address_task_ready),
    .io_read_address_task_valid(argRouteServers_0_io_read_address_task_valid),
    .io_read_address_task_bits(argRouteServers_0_io_read_address_task_bits),
    .io_read_data_task_ready(argRouteServers_0_io_read_data_task_ready),
    .io_read_data_task_valid(argRouteServers_0_io_read_data_task_valid),
    .io_read_data_task_bits(argRouteServers_0_io_read_data_task_bits)
  );
  argRouteVirtServerV2 argRouteServers_1 ( // @[syncSide.scala 55:15]
    .clock(argRouteServers_1_clock),
    .reset(argRouteServers_1_reset),
    .io_connNetwork_ready(argRouteServers_1_io_connNetwork_ready),
    .io_connNetwork_valid(argRouteServers_1_io_connNetwork_valid),
    .io_connNetwork_bits(argRouteServers_1_io_connNetwork_bits),
    .io_connStealNtw_ctrl_serveStealReq_ready(argRouteServers_1_io_connStealNtw_ctrl_serveStealReq_ready),
    .io_connStealNtw_ctrl_serveStealReq_valid(argRouteServers_1_io_connStealNtw_ctrl_serveStealReq_valid),
    .io_connStealNtw_data_qOutTask_ready(argRouteServers_1_io_connStealNtw_data_qOutTask_ready),
    .io_connStealNtw_data_qOutTask_valid(argRouteServers_1_io_connStealNtw_data_qOutTask_valid),
    .io_connStealNtw_data_qOutTask_bits(argRouteServers_1_io_connStealNtw_data_qOutTask_bits),
    .io_read_address_ready(argRouteServers_1_io_read_address_ready),
    .io_read_address_valid(argRouteServers_1_io_read_address_valid),
    .io_read_address_bits(argRouteServers_1_io_read_address_bits),
    .io_read_data_ready(argRouteServers_1_io_read_data_ready),
    .io_read_data_valid(argRouteServers_1_io_read_data_valid),
    .io_read_data_bits(argRouteServers_1_io_read_data_bits),
    .io_write_address_ready(argRouteServers_1_io_write_address_ready),
    .io_write_address_valid(argRouteServers_1_io_write_address_valid),
    .io_write_address_bits(argRouteServers_1_io_write_address_bits),
    .io_write_data_ready(argRouteServers_1_io_write_data_ready),
    .io_write_data_valid(argRouteServers_1_io_write_data_valid),
    .io_write_data_bits(argRouteServers_1_io_write_data_bits),
    .io_read_address_task_ready(argRouteServers_1_io_read_address_task_ready),
    .io_read_address_task_valid(argRouteServers_1_io_read_address_task_valid),
    .io_read_address_task_bits(argRouteServers_1_io_read_address_task_bits),
    .io_read_data_task_ready(argRouteServers_1_io_read_data_task_ready),
    .io_read_data_task_valid(argRouteServers_1_io_read_data_task_valid),
    .io_read_data_task_bits(argRouteServers_1_io_read_data_task_bits)
  );
  readyValidMem_2 argRouteRvm_0 ( // @[syncSide.scala 65:67]
    .clock(argRouteRvm_0_clock),
    .reset(argRouteRvm_0_reset),
    .io_read_address_ready(argRouteRvm_0_io_read_address_ready),
    .io_read_address_valid(argRouteRvm_0_io_read_address_valid),
    .io_read_address_bits(argRouteRvm_0_io_read_address_bits),
    .io_read_data_ready(argRouteRvm_0_io_read_data_ready),
    .io_read_data_valid(argRouteRvm_0_io_read_data_valid),
    .io_read_data_bits(argRouteRvm_0_io_read_data_bits),
    .io_write_address_ready(argRouteRvm_0_io_write_address_ready),
    .io_write_address_valid(argRouteRvm_0_io_write_address_valid),
    .io_write_address_bits(argRouteRvm_0_io_write_address_bits),
    .io_write_data_ready(argRouteRvm_0_io_write_data_ready),
    .io_write_data_valid(argRouteRvm_0_io_write_data_valid),
    .io_write_data_bits(argRouteRvm_0_io_write_data_bits),
    .axi_ARREADY(argRouteRvm_0_axi_ARREADY),
    .axi_ARVALID(argRouteRvm_0_axi_ARVALID),
    .axi_ARADDR(argRouteRvm_0_axi_ARADDR),
    .axi_RREADY(argRouteRvm_0_axi_RREADY),
    .axi_RVALID(argRouteRvm_0_axi_RVALID),
    .axi_RDATA(argRouteRvm_0_axi_RDATA),
    .axi_AWREADY(argRouteRvm_0_axi_AWREADY),
    .axi_AWVALID(argRouteRvm_0_axi_AWVALID),
    .axi_AWADDR(argRouteRvm_0_axi_AWADDR),
    .axi_WREADY(argRouteRvm_0_axi_WREADY),
    .axi_WVALID(argRouteRvm_0_axi_WVALID),
    .axi_WDATA(argRouteRvm_0_axi_WDATA),
    .axi_BVALID(argRouteRvm_0_axi_BVALID)
  );
  readyValidMem_2 argRouteRvm_1 ( // @[syncSide.scala 65:67]
    .clock(argRouteRvm_1_clock),
    .reset(argRouteRvm_1_reset),
    .io_read_address_ready(argRouteRvm_1_io_read_address_ready),
    .io_read_address_valid(argRouteRvm_1_io_read_address_valid),
    .io_read_address_bits(argRouteRvm_1_io_read_address_bits),
    .io_read_data_ready(argRouteRvm_1_io_read_data_ready),
    .io_read_data_valid(argRouteRvm_1_io_read_data_valid),
    .io_read_data_bits(argRouteRvm_1_io_read_data_bits),
    .io_write_address_ready(argRouteRvm_1_io_write_address_ready),
    .io_write_address_valid(argRouteRvm_1_io_write_address_valid),
    .io_write_address_bits(argRouteRvm_1_io_write_address_bits),
    .io_write_data_ready(argRouteRvm_1_io_write_data_ready),
    .io_write_data_valid(argRouteRvm_1_io_write_data_valid),
    .io_write_data_bits(argRouteRvm_1_io_write_data_bits),
    .axi_ARREADY(argRouteRvm_1_axi_ARREADY),
    .axi_ARVALID(argRouteRvm_1_axi_ARVALID),
    .axi_ARADDR(argRouteRvm_1_axi_ARADDR),
    .axi_RREADY(argRouteRvm_1_axi_RREADY),
    .axi_RVALID(argRouteRvm_1_axi_RVALID),
    .axi_RDATA(argRouteRvm_1_axi_RDATA),
    .axi_AWREADY(argRouteRvm_1_axi_AWREADY),
    .axi_AWVALID(argRouteRvm_1_axi_AWVALID),
    .axi_AWADDR(argRouteRvm_1_axi_AWADDR),
    .axi_WREADY(argRouteRvm_1_axi_WREADY),
    .axi_WVALID(argRouteRvm_1_axi_WVALID),
    .axi_WDATA(argRouteRvm_1_axi_WDATA),
    .axi_BVALID(argRouteRvm_1_axi_BVALID)
  );
  readyValidMem_4 argRouteRvmReadOnly_0 ( // @[syncSide.scala 66:69]
    .io_read_address_ready(argRouteRvmReadOnly_0_io_read_address_ready),
    .io_read_address_valid(argRouteRvmReadOnly_0_io_read_address_valid),
    .io_read_address_bits(argRouteRvmReadOnly_0_io_read_address_bits),
    .io_read_data_ready(argRouteRvmReadOnly_0_io_read_data_ready),
    .io_read_data_valid(argRouteRvmReadOnly_0_io_read_data_valid),
    .io_read_data_bits(argRouteRvmReadOnly_0_io_read_data_bits),
    .axi_ARREADY(argRouteRvmReadOnly_0_axi_ARREADY),
    .axi_ARVALID(argRouteRvmReadOnly_0_axi_ARVALID),
    .axi_ARADDR(argRouteRvmReadOnly_0_axi_ARADDR),
    .axi_RREADY(argRouteRvmReadOnly_0_axi_RREADY),
    .axi_RVALID(argRouteRvmReadOnly_0_axi_RVALID),
    .axi_RDATA(argRouteRvmReadOnly_0_axi_RDATA)
  );
  readyValidMem_4 argRouteRvmReadOnly_1 ( // @[syncSide.scala 66:69]
    .io_read_address_ready(argRouteRvmReadOnly_1_io_read_address_ready),
    .io_read_address_valid(argRouteRvmReadOnly_1_io_read_address_valid),
    .io_read_address_bits(argRouteRvmReadOnly_1_io_read_address_bits),
    .io_read_data_ready(argRouteRvmReadOnly_1_io_read_data_ready),
    .io_read_data_valid(argRouteRvmReadOnly_1_io_read_data_valid),
    .io_read_data_bits(argRouteRvmReadOnly_1_io_read_data_bits),
    .axi_ARREADY(argRouteRvmReadOnly_1_axi_ARREADY),
    .axi_ARVALID(argRouteRvmReadOnly_1_axi_ARVALID),
    .axi_ARADDR(argRouteRvmReadOnly_1_axi_ARADDR),
    .axi_RREADY(argRouteRvmReadOnly_1_axi_RREADY),
    .axi_RVALID(argRouteRvmReadOnly_1_axi_RVALID),
    .axi_RDATA(argRouteRvmReadOnly_1_axi_RDATA)
  );
  assign io_addrIn_0_TREADY = argSide_io_connPE_0_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_1_TREADY = argSide_io_connPE_1_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_2_TREADY = argSide_io_connPE_2_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_3_TREADY = argSide_io_connPE_3_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_4_TREADY = argSide_io_connPE_4_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_5_TREADY = argSide_io_connPE_5_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_6_TREADY = argSide_io_connPE_6_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_7_TREADY = argSide_io_connPE_7_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_8_TREADY = argSide_io_connPE_8_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_9_TREADY = argSide_io_connPE_9_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_10_TREADY = argSide_io_connPE_10_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_11_TREADY = argSide_io_connPE_11_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_12_TREADY = argSide_io_connPE_12_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_13_TREADY = argSide_io_connPE_13_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_14_TREADY = argSide_io_connPE_14_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_15_TREADY = argSide_io_connPE_15_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_16_TREADY = argSide_io_connPE_16_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_17_TREADY = argSide_io_connPE_17_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_18_TREADY = argSide_io_connPE_18_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_19_TREADY = argSide_io_connPE_19_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_20_TREADY = argSide_io_connPE_20_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_21_TREADY = argSide_io_connPE_21_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_22_TREADY = argSide_io_connPE_22_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_23_TREADY = argSide_io_connPE_23_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_24_TREADY = argSide_io_connPE_24_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_25_TREADY = argSide_io_connPE_25_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_26_TREADY = argSide_io_connPE_26_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_27_TREADY = argSide_io_connPE_27_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_28_TREADY = argSide_io_connPE_28_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_29_TREADY = argSide_io_connPE_29_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_30_TREADY = argSide_io_connPE_30_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_31_TREADY = argSide_io_connPE_31_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_32_TREADY = argSide_io_connPE_32_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_33_TREADY = argSide_io_connPE_33_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_34_TREADY = argSide_io_connPE_34_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_35_TREADY = argSide_io_connPE_35_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_36_TREADY = argSide_io_connPE_36_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_37_TREADY = argSide_io_connPE_37_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_38_TREADY = argSide_io_connPE_38_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_39_TREADY = argSide_io_connPE_39_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_40_TREADY = argSide_io_connPE_40_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_41_TREADY = argSide_io_connPE_41_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_42_TREADY = argSide_io_connPE_42_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_43_TREADY = argSide_io_connPE_43_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_44_TREADY = argSide_io_connPE_44_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_45_TREADY = argSide_io_connPE_45_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_46_TREADY = argSide_io_connPE_46_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_47_TREADY = argSide_io_connPE_47_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_48_TREADY = argSide_io_connPE_48_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_49_TREADY = argSide_io_connPE_49_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_50_TREADY = argSide_io_connPE_50_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_51_TREADY = argSide_io_connPE_51_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_52_TREADY = argSide_io_connPE_52_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_53_TREADY = argSide_io_connPE_53_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_54_TREADY = argSide_io_connPE_54_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_55_TREADY = argSide_io_connPE_55_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_56_TREADY = argSide_io_connPE_56_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_57_TREADY = argSide_io_connPE_57_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_58_TREADY = argSide_io_connPE_58_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_59_TREADY = argSide_io_connPE_59_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_60_TREADY = argSide_io_connPE_60_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_61_TREADY = argSide_io_connPE_61_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_62_TREADY = argSide_io_connPE_62_ready; // @[syncSide.scala 83:30]
  assign io_addrIn_63_TREADY = argSide_io_connPE_63_ready; // @[syncSide.scala 83:30]
  assign io_axi_full_argRoute_0_ARVALID = argRouteRvm_0_axi_ARVALID; // @[syncSide.scala 69:45]
  assign io_axi_full_argRoute_0_ARADDR = argRouteRvm_0_axi_ARADDR; // @[syncSide.scala 69:45]
  assign io_axi_full_argRoute_0_RREADY = argRouteRvm_0_axi_RREADY; // @[syncSide.scala 69:45]
  assign io_axi_full_argRoute_0_AWVALID = argRouteRvm_0_axi_AWVALID; // @[syncSide.scala 69:45]
  assign io_axi_full_argRoute_0_AWADDR = argRouteRvm_0_axi_AWADDR; // @[syncSide.scala 69:45]
  assign io_axi_full_argRoute_0_WVALID = argRouteRvm_0_axi_WVALID; // @[syncSide.scala 69:45]
  assign io_axi_full_argRoute_0_WDATA = argRouteRvm_0_axi_WDATA; // @[syncSide.scala 69:45]
  assign io_axi_full_argRoute_1_ARVALID = argRouteRvm_1_axi_ARVALID; // @[syncSide.scala 69:45]
  assign io_axi_full_argRoute_1_ARADDR = argRouteRvm_1_axi_ARADDR; // @[syncSide.scala 69:45]
  assign io_axi_full_argRoute_1_RREADY = argRouteRvm_1_axi_RREADY; // @[syncSide.scala 69:45]
  assign io_axi_full_argRoute_1_AWVALID = argRouteRvm_1_axi_AWVALID; // @[syncSide.scala 69:45]
  assign io_axi_full_argRoute_1_AWADDR = argRouteRvm_1_axi_AWADDR; // @[syncSide.scala 69:45]
  assign io_axi_full_argRoute_1_WVALID = argRouteRvm_1_axi_WVALID; // @[syncSide.scala 69:45]
  assign io_axi_full_argRoute_1_WDATA = argRouteRvm_1_axi_WDATA; // @[syncSide.scala 69:45]
  assign io_axi_full_argRoute_2_ARVALID = argRouteRvmReadOnly_0_axi_ARVALID; // @[syncSide.scala 77:55]
  assign io_axi_full_argRoute_2_ARADDR = argRouteRvmReadOnly_0_axi_ARADDR; // @[syncSide.scala 77:55]
  assign io_axi_full_argRoute_2_RREADY = argRouteRvmReadOnly_0_axi_RREADY; // @[syncSide.scala 77:55]
  assign io_axi_full_argRoute_3_ARVALID = argRouteRvmReadOnly_1_axi_ARVALID; // @[syncSide.scala 77:55]
  assign io_axi_full_argRoute_3_ARADDR = argRouteRvmReadOnly_1_axi_ARADDR; // @[syncSide.scala 77:55]
  assign io_axi_full_argRoute_3_RREADY = argRouteRvmReadOnly_1_axi_RREADY; // @[syncSide.scala 77:55]
  assign connStealNtw_0_ctrl_serveStealReq_valid = argRouteServers_0_io_connStealNtw_ctrl_serveStealReq_valid; // @[syncSide.scala 75:45]
  assign connStealNtw_0_data_qOutTask_valid = argRouteServers_0_io_connStealNtw_data_qOutTask_valid; // @[syncSide.scala 75:45]
  assign connStealNtw_0_data_qOutTask_bits = argRouteServers_0_io_connStealNtw_data_qOutTask_bits; // @[syncSide.scala 75:45]
  assign connStealNtw_1_ctrl_serveStealReq_valid = argRouteServers_1_io_connStealNtw_ctrl_serveStealReq_valid; // @[syncSide.scala 75:45]
  assign connStealNtw_1_data_qOutTask_valid = argRouteServers_1_io_connStealNtw_data_qOutTask_valid; // @[syncSide.scala 75:45]
  assign connStealNtw_1_data_qOutTask_bits = argRouteServers_1_io_connStealNtw_data_qOutTask_bits; // @[syncSide.scala 75:45]
  assign argSide_clock = clock;
  assign argSide_reset = reset;
  assign argSide_io_connVAS_0_ready = argRouteServers_0_io_connNetwork_ready; // @[syncSide.scala 74:45]
  assign argSide_io_connVAS_1_ready = argRouteServers_1_io_connNetwork_ready; // @[syncSide.scala 74:45]
  assign argSide_io_connPE_0_valid = io_addrIn_0_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_0_bits = io_addrIn_0_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_1_valid = io_addrIn_1_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_1_bits = io_addrIn_1_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_2_valid = io_addrIn_2_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_2_bits = io_addrIn_2_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_3_valid = io_addrIn_3_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_3_bits = io_addrIn_3_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_4_valid = io_addrIn_4_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_4_bits = io_addrIn_4_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_5_valid = io_addrIn_5_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_5_bits = io_addrIn_5_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_6_valid = io_addrIn_6_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_6_bits = io_addrIn_6_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_7_valid = io_addrIn_7_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_7_bits = io_addrIn_7_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_8_valid = io_addrIn_8_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_8_bits = io_addrIn_8_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_9_valid = io_addrIn_9_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_9_bits = io_addrIn_9_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_10_valid = io_addrIn_10_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_10_bits = io_addrIn_10_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_11_valid = io_addrIn_11_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_11_bits = io_addrIn_11_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_12_valid = io_addrIn_12_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_12_bits = io_addrIn_12_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_13_valid = io_addrIn_13_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_13_bits = io_addrIn_13_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_14_valid = io_addrIn_14_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_14_bits = io_addrIn_14_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_15_valid = io_addrIn_15_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_15_bits = io_addrIn_15_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_16_valid = io_addrIn_16_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_16_bits = io_addrIn_16_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_17_valid = io_addrIn_17_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_17_bits = io_addrIn_17_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_18_valid = io_addrIn_18_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_18_bits = io_addrIn_18_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_19_valid = io_addrIn_19_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_19_bits = io_addrIn_19_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_20_valid = io_addrIn_20_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_20_bits = io_addrIn_20_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_21_valid = io_addrIn_21_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_21_bits = io_addrIn_21_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_22_valid = io_addrIn_22_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_22_bits = io_addrIn_22_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_23_valid = io_addrIn_23_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_23_bits = io_addrIn_23_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_24_valid = io_addrIn_24_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_24_bits = io_addrIn_24_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_25_valid = io_addrIn_25_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_25_bits = io_addrIn_25_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_26_valid = io_addrIn_26_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_26_bits = io_addrIn_26_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_27_valid = io_addrIn_27_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_27_bits = io_addrIn_27_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_28_valid = io_addrIn_28_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_28_bits = io_addrIn_28_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_29_valid = io_addrIn_29_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_29_bits = io_addrIn_29_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_30_valid = io_addrIn_30_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_30_bits = io_addrIn_30_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_31_valid = io_addrIn_31_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_31_bits = io_addrIn_31_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_32_valid = io_addrIn_32_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_32_bits = io_addrIn_32_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_33_valid = io_addrIn_33_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_33_bits = io_addrIn_33_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_34_valid = io_addrIn_34_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_34_bits = io_addrIn_34_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_35_valid = io_addrIn_35_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_35_bits = io_addrIn_35_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_36_valid = io_addrIn_36_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_36_bits = io_addrIn_36_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_37_valid = io_addrIn_37_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_37_bits = io_addrIn_37_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_38_valid = io_addrIn_38_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_38_bits = io_addrIn_38_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_39_valid = io_addrIn_39_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_39_bits = io_addrIn_39_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_40_valid = io_addrIn_40_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_40_bits = io_addrIn_40_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_41_valid = io_addrIn_41_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_41_bits = io_addrIn_41_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_42_valid = io_addrIn_42_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_42_bits = io_addrIn_42_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_43_valid = io_addrIn_43_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_43_bits = io_addrIn_43_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_44_valid = io_addrIn_44_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_44_bits = io_addrIn_44_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_45_valid = io_addrIn_45_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_45_bits = io_addrIn_45_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_46_valid = io_addrIn_46_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_46_bits = io_addrIn_46_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_47_valid = io_addrIn_47_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_47_bits = io_addrIn_47_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_48_valid = io_addrIn_48_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_48_bits = io_addrIn_48_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_49_valid = io_addrIn_49_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_49_bits = io_addrIn_49_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_50_valid = io_addrIn_50_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_50_bits = io_addrIn_50_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_51_valid = io_addrIn_51_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_51_bits = io_addrIn_51_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_52_valid = io_addrIn_52_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_52_bits = io_addrIn_52_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_53_valid = io_addrIn_53_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_53_bits = io_addrIn_53_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_54_valid = io_addrIn_54_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_54_bits = io_addrIn_54_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_55_valid = io_addrIn_55_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_55_bits = io_addrIn_55_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_56_valid = io_addrIn_56_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_56_bits = io_addrIn_56_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_57_valid = io_addrIn_57_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_57_bits = io_addrIn_57_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_58_valid = io_addrIn_58_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_58_bits = io_addrIn_58_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_59_valid = io_addrIn_59_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_59_bits = io_addrIn_59_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_60_valid = io_addrIn_60_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_60_bits = io_addrIn_60_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_61_valid = io_addrIn_61_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_61_bits = io_addrIn_61_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_62_valid = io_addrIn_62_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_62_bits = io_addrIn_62_TDATA; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_63_valid = io_addrIn_63_TVALID; // @[syncSide.scala 83:30]
  assign argSide_io_connPE_63_bits = io_addrIn_63_TDATA; // @[syncSide.scala 83:30]
  assign argRouteServers_0_clock = clock;
  assign argRouteServers_0_reset = reset;
  assign argRouteServers_0_io_connNetwork_valid = argSide_io_connVAS_0_valid; // @[syncSide.scala 74:45]
  assign argRouteServers_0_io_connNetwork_bits = argSide_io_connVAS_0_bits; // @[syncSide.scala 74:45]
  assign argRouteServers_0_io_connStealNtw_ctrl_serveStealReq_ready = connStealNtw_0_ctrl_serveStealReq_ready; // @[syncSide.scala 75:45]
  assign argRouteServers_0_io_connStealNtw_data_qOutTask_ready = connStealNtw_0_data_qOutTask_ready; // @[syncSide.scala 75:45]
  assign argRouteServers_0_io_read_address_ready = argRouteRvm_0_io_read_address_ready; // @[syncSide.scala 70:45]
  assign argRouteServers_0_io_read_data_valid = argRouteRvm_0_io_read_data_valid; // @[syncSide.scala 71:45]
  assign argRouteServers_0_io_read_data_bits = argRouteRvm_0_io_read_data_bits; // @[syncSide.scala 71:45]
  assign argRouteServers_0_io_write_address_ready = argRouteRvm_0_io_write_address_ready; // @[syncSide.scala 72:45]
  assign argRouteServers_0_io_write_data_ready = argRouteRvm_0_io_write_data_ready; // @[syncSide.scala 73:45]
  assign argRouteServers_0_io_read_address_task_ready = argRouteRvmReadOnly_0_io_read_address_ready; // @[syncSide.scala 78:53]
  assign argRouteServers_0_io_read_data_task_valid = argRouteRvmReadOnly_0_io_read_data_valid; // @[syncSide.scala 79:53]
  assign argRouteServers_0_io_read_data_task_bits = argRouteRvmReadOnly_0_io_read_data_bits; // @[syncSide.scala 79:53]
  assign argRouteServers_1_clock = clock;
  assign argRouteServers_1_reset = reset;
  assign argRouteServers_1_io_connNetwork_valid = argSide_io_connVAS_1_valid; // @[syncSide.scala 74:45]
  assign argRouteServers_1_io_connNetwork_bits = argSide_io_connVAS_1_bits; // @[syncSide.scala 74:45]
  assign argRouteServers_1_io_connStealNtw_ctrl_serveStealReq_ready = connStealNtw_1_ctrl_serveStealReq_ready; // @[syncSide.scala 75:45]
  assign argRouteServers_1_io_connStealNtw_data_qOutTask_ready = connStealNtw_1_data_qOutTask_ready; // @[syncSide.scala 75:45]
  assign argRouteServers_1_io_read_address_ready = argRouteRvm_1_io_read_address_ready; // @[syncSide.scala 70:45]
  assign argRouteServers_1_io_read_data_valid = argRouteRvm_1_io_read_data_valid; // @[syncSide.scala 71:45]
  assign argRouteServers_1_io_read_data_bits = argRouteRvm_1_io_read_data_bits; // @[syncSide.scala 71:45]
  assign argRouteServers_1_io_write_address_ready = argRouteRvm_1_io_write_address_ready; // @[syncSide.scala 72:45]
  assign argRouteServers_1_io_write_data_ready = argRouteRvm_1_io_write_data_ready; // @[syncSide.scala 73:45]
  assign argRouteServers_1_io_read_address_task_ready = argRouteRvmReadOnly_1_io_read_address_ready; // @[syncSide.scala 78:53]
  assign argRouteServers_1_io_read_data_task_valid = argRouteRvmReadOnly_1_io_read_data_valid; // @[syncSide.scala 79:53]
  assign argRouteServers_1_io_read_data_task_bits = argRouteRvmReadOnly_1_io_read_data_bits; // @[syncSide.scala 79:53]
  assign argRouteRvm_0_clock = clock;
  assign argRouteRvm_0_reset = reset;
  assign argRouteRvm_0_io_read_address_valid = argRouteServers_0_io_read_address_valid; // @[syncSide.scala 70:45]
  assign argRouteRvm_0_io_read_address_bits = argRouteServers_0_io_read_address_bits; // @[syncSide.scala 70:45]
  assign argRouteRvm_0_io_read_data_ready = argRouteServers_0_io_read_data_ready; // @[syncSide.scala 71:45]
  assign argRouteRvm_0_io_write_address_valid = argRouteServers_0_io_write_address_valid; // @[syncSide.scala 72:45]
  assign argRouteRvm_0_io_write_address_bits = argRouteServers_0_io_write_address_bits; // @[syncSide.scala 72:45]
  assign argRouteRvm_0_io_write_data_valid = argRouteServers_0_io_write_data_valid; // @[syncSide.scala 73:45]
  assign argRouteRvm_0_io_write_data_bits = argRouteServers_0_io_write_data_bits; // @[syncSide.scala 73:45]
  assign argRouteRvm_0_axi_ARREADY = io_axi_full_argRoute_0_ARREADY; // @[syncSide.scala 69:45]
  assign argRouteRvm_0_axi_RVALID = io_axi_full_argRoute_0_RVALID; // @[syncSide.scala 69:45]
  assign argRouteRvm_0_axi_RDATA = io_axi_full_argRoute_0_RDATA; // @[syncSide.scala 69:45]
  assign argRouteRvm_0_axi_AWREADY = io_axi_full_argRoute_0_AWREADY; // @[syncSide.scala 69:45]
  assign argRouteRvm_0_axi_WREADY = io_axi_full_argRoute_0_WREADY; // @[syncSide.scala 69:45]
  assign argRouteRvm_0_axi_BVALID = io_axi_full_argRoute_0_BVALID; // @[syncSide.scala 69:45]
  assign argRouteRvm_1_clock = clock;
  assign argRouteRvm_1_reset = reset;
  assign argRouteRvm_1_io_read_address_valid = argRouteServers_1_io_read_address_valid; // @[syncSide.scala 70:45]
  assign argRouteRvm_1_io_read_address_bits = argRouteServers_1_io_read_address_bits; // @[syncSide.scala 70:45]
  assign argRouteRvm_1_io_read_data_ready = argRouteServers_1_io_read_data_ready; // @[syncSide.scala 71:45]
  assign argRouteRvm_1_io_write_address_valid = argRouteServers_1_io_write_address_valid; // @[syncSide.scala 72:45]
  assign argRouteRvm_1_io_write_address_bits = argRouteServers_1_io_write_address_bits; // @[syncSide.scala 72:45]
  assign argRouteRvm_1_io_write_data_valid = argRouteServers_1_io_write_data_valid; // @[syncSide.scala 73:45]
  assign argRouteRvm_1_io_write_data_bits = argRouteServers_1_io_write_data_bits; // @[syncSide.scala 73:45]
  assign argRouteRvm_1_axi_ARREADY = io_axi_full_argRoute_1_ARREADY; // @[syncSide.scala 69:45]
  assign argRouteRvm_1_axi_RVALID = io_axi_full_argRoute_1_RVALID; // @[syncSide.scala 69:45]
  assign argRouteRvm_1_axi_RDATA = io_axi_full_argRoute_1_RDATA; // @[syncSide.scala 69:45]
  assign argRouteRvm_1_axi_AWREADY = io_axi_full_argRoute_1_AWREADY; // @[syncSide.scala 69:45]
  assign argRouteRvm_1_axi_WREADY = io_axi_full_argRoute_1_WREADY; // @[syncSide.scala 69:45]
  assign argRouteRvm_1_axi_BVALID = io_axi_full_argRoute_1_BVALID; // @[syncSide.scala 69:45]
  assign argRouteRvmReadOnly_0_io_read_address_valid = argRouteServers_0_io_read_address_task_valid; // @[syncSide.scala 78:53]
  assign argRouteRvmReadOnly_0_io_read_address_bits = argRouteServers_0_io_read_address_task_bits; // @[syncSide.scala 78:53]
  assign argRouteRvmReadOnly_0_io_read_data_ready = argRouteServers_0_io_read_data_task_ready; // @[syncSide.scala 79:53]
  assign argRouteRvmReadOnly_0_axi_ARREADY = io_axi_full_argRoute_2_ARREADY; // @[syncSide.scala 77:55]
  assign argRouteRvmReadOnly_0_axi_RVALID = io_axi_full_argRoute_2_RVALID; // @[syncSide.scala 77:55]
  assign argRouteRvmReadOnly_0_axi_RDATA = io_axi_full_argRoute_2_RDATA; // @[syncSide.scala 77:55]
  assign argRouteRvmReadOnly_1_io_read_address_valid = argRouteServers_1_io_read_address_task_valid; // @[syncSide.scala 78:53]
  assign argRouteRvmReadOnly_1_io_read_address_bits = argRouteServers_1_io_read_address_task_bits; // @[syncSide.scala 78:53]
  assign argRouteRvmReadOnly_1_io_read_data_ready = argRouteServers_1_io_read_data_task_ready; // @[syncSide.scala 79:53]
  assign argRouteRvmReadOnly_1_axi_ARREADY = io_axi_full_argRoute_3_ARREADY; // @[syncSide.scala 77:55]
  assign argRouteRvmReadOnly_1_axi_RVALID = io_axi_full_argRoute_3_RVALID; // @[syncSide.scala 77:55]
  assign argRouteRvmReadOnly_1_axi_RDATA = io_axi_full_argRoute_3_RDATA; // @[syncSide.scala 77:55]
endmodule
module fullSysGen(
  input          clock,
  input          reset,
  output         task_stealSide_axi_mgmt_vss_0_ARREADY,
  input          task_stealSide_axi_mgmt_vss_0_ARVALID,
  input  [5:0]   task_stealSide_axi_mgmt_vss_0_ARADDR,
  input  [2:0]   task_stealSide_axi_mgmt_vss_0_ARPROT,
  input          task_stealSide_axi_mgmt_vss_0_RREADY,
  output         task_stealSide_axi_mgmt_vss_0_RVALID,
  output [63:0]  task_stealSide_axi_mgmt_vss_0_RDATA,
  output [1:0]   task_stealSide_axi_mgmt_vss_0_RRESP,
  output         task_stealSide_axi_mgmt_vss_0_AWREADY,
  input          task_stealSide_axi_mgmt_vss_0_AWVALID,
  input  [5:0]   task_stealSide_axi_mgmt_vss_0_AWADDR,
  input  [2:0]   task_stealSide_axi_mgmt_vss_0_AWPROT,
  output         task_stealSide_axi_mgmt_vss_0_WREADY,
  input          task_stealSide_axi_mgmt_vss_0_WVALID,
  input  [63:0]  task_stealSide_axi_mgmt_vss_0_WDATA,
  input  [7:0]   task_stealSide_axi_mgmt_vss_0_WSTRB,
  input          task_stealSide_axi_mgmt_vss_0_BREADY,
  output         task_stealSide_axi_mgmt_vss_0_BVALID,
  output [1:0]   task_stealSide_axi_mgmt_vss_0_BRESP,
  input          task_stealSide_vss_axi_full_0_ARREADY,
  output         task_stealSide_vss_axi_full_0_ARVALID,
  output [3:0]   task_stealSide_vss_axi_full_0_ARID,
  output [63:0]  task_stealSide_vss_axi_full_0_ARADDR,
  output [7:0]   task_stealSide_vss_axi_full_0_ARLEN,
  output [2:0]   task_stealSide_vss_axi_full_0_ARSIZE,
  output [1:0]   task_stealSide_vss_axi_full_0_ARBURST,
  output         task_stealSide_vss_axi_full_0_ARLOCK,
  output [3:0]   task_stealSide_vss_axi_full_0_ARCACHE,
  output [2:0]   task_stealSide_vss_axi_full_0_ARPROT,
  output [3:0]   task_stealSide_vss_axi_full_0_ARQOS,
  output [3:0]   task_stealSide_vss_axi_full_0_ARREGION,
  output         task_stealSide_vss_axi_full_0_RREADY,
  input          task_stealSide_vss_axi_full_0_RVALID,
  input  [3:0]   task_stealSide_vss_axi_full_0_RID,
  input  [255:0] task_stealSide_vss_axi_full_0_RDATA,
  input  [1:0]   task_stealSide_vss_axi_full_0_RRESP,
  input          task_stealSide_vss_axi_full_0_RLAST,
  input          task_stealSide_vss_axi_full_0_AWREADY,
  output         task_stealSide_vss_axi_full_0_AWVALID,
  output [3:0]   task_stealSide_vss_axi_full_0_AWID,
  output [63:0]  task_stealSide_vss_axi_full_0_AWADDR,
  output [7:0]   task_stealSide_vss_axi_full_0_AWLEN,
  output [2:0]   task_stealSide_vss_axi_full_0_AWSIZE,
  output [1:0]   task_stealSide_vss_axi_full_0_AWBURST,
  output         task_stealSide_vss_axi_full_0_AWLOCK,
  output [3:0]   task_stealSide_vss_axi_full_0_AWCACHE,
  output [2:0]   task_stealSide_vss_axi_full_0_AWPROT,
  output [3:0]   task_stealSide_vss_axi_full_0_AWQOS,
  output [3:0]   task_stealSide_vss_axi_full_0_AWREGION,
  input          task_stealSide_vss_axi_full_0_WREADY,
  output         task_stealSide_vss_axi_full_0_WVALID,
  output [3:0]   task_stealSide_vss_axi_full_0_WID,
  output [255:0] task_stealSide_vss_axi_full_0_WDATA,
  output [31:0]  task_stealSide_vss_axi_full_0_WSTRB,
  output         task_stealSide_vss_axi_full_0_WLAST,
  output         task_stealSide_vss_axi_full_0_BREADY,
  input          task_stealSide_vss_axi_full_0_BVALID,
  input  [3:0]   task_stealSide_vss_axi_full_0_BID,
  input  [1:0]   task_stealSide_vss_axi_full_0_BRESP,
  input          task_stealSide_taskOut_0_TREADY,
  output         task_stealSide_taskOut_0_TVALID,
  output [255:0] task_stealSide_taskOut_0_TDATA,
  input          task_stealSide_taskOut_1_TREADY,
  output         task_stealSide_taskOut_1_TVALID,
  output [255:0] task_stealSide_taskOut_1_TDATA,
  input          task_stealSide_taskOut_2_TREADY,
  output         task_stealSide_taskOut_2_TVALID,
  output [255:0] task_stealSide_taskOut_2_TDATA,
  input          task_stealSide_taskOut_3_TREADY,
  output         task_stealSide_taskOut_3_TVALID,
  output [255:0] task_stealSide_taskOut_3_TDATA,
  input          task_stealSide_taskOut_4_TREADY,
  output         task_stealSide_taskOut_4_TVALID,
  output [255:0] task_stealSide_taskOut_4_TDATA,
  input          task_stealSide_taskOut_5_TREADY,
  output         task_stealSide_taskOut_5_TVALID,
  output [255:0] task_stealSide_taskOut_5_TDATA,
  input          task_stealSide_taskOut_6_TREADY,
  output         task_stealSide_taskOut_6_TVALID,
  output [255:0] task_stealSide_taskOut_6_TDATA,
  input          task_stealSide_taskOut_7_TREADY,
  output         task_stealSide_taskOut_7_TVALID,
  output [255:0] task_stealSide_taskOut_7_TDATA,
  input          task_stealSide_taskOut_8_TREADY,
  output         task_stealSide_taskOut_8_TVALID,
  output [255:0] task_stealSide_taskOut_8_TDATA,
  input          task_stealSide_taskOut_9_TREADY,
  output         task_stealSide_taskOut_9_TVALID,
  output [255:0] task_stealSide_taskOut_9_TDATA,
  input          task_stealSide_taskOut_10_TREADY,
  output         task_stealSide_taskOut_10_TVALID,
  output [255:0] task_stealSide_taskOut_10_TDATA,
  input          task_stealSide_taskOut_11_TREADY,
  output         task_stealSide_taskOut_11_TVALID,
  output [255:0] task_stealSide_taskOut_11_TDATA,
  input          task_stealSide_taskOut_12_TREADY,
  output         task_stealSide_taskOut_12_TVALID,
  output [255:0] task_stealSide_taskOut_12_TDATA,
  input          task_stealSide_taskOut_13_TREADY,
  output         task_stealSide_taskOut_13_TVALID,
  output [255:0] task_stealSide_taskOut_13_TDATA,
  input          task_stealSide_taskOut_14_TREADY,
  output         task_stealSide_taskOut_14_TVALID,
  output [255:0] task_stealSide_taskOut_14_TDATA,
  input          task_stealSide_taskOut_15_TREADY,
  output         task_stealSide_taskOut_15_TVALID,
  output [255:0] task_stealSide_taskOut_15_TDATA,
  input          task_stealSide_taskOut_16_TREADY,
  output         task_stealSide_taskOut_16_TVALID,
  output [255:0] task_stealSide_taskOut_16_TDATA,
  input          task_stealSide_taskOut_17_TREADY,
  output         task_stealSide_taskOut_17_TVALID,
  output [255:0] task_stealSide_taskOut_17_TDATA,
  input          task_stealSide_taskOut_18_TREADY,
  output         task_stealSide_taskOut_18_TVALID,
  output [255:0] task_stealSide_taskOut_18_TDATA,
  input          task_stealSide_taskOut_19_TREADY,
  output         task_stealSide_taskOut_19_TVALID,
  output [255:0] task_stealSide_taskOut_19_TDATA,
  input          task_stealSide_taskOut_20_TREADY,
  output         task_stealSide_taskOut_20_TVALID,
  output [255:0] task_stealSide_taskOut_20_TDATA,
  input          task_stealSide_taskOut_21_TREADY,
  output         task_stealSide_taskOut_21_TVALID,
  output [255:0] task_stealSide_taskOut_21_TDATA,
  input          task_stealSide_taskOut_22_TREADY,
  output         task_stealSide_taskOut_22_TVALID,
  output [255:0] task_stealSide_taskOut_22_TDATA,
  input          task_stealSide_taskOut_23_TREADY,
  output         task_stealSide_taskOut_23_TVALID,
  output [255:0] task_stealSide_taskOut_23_TDATA,
  input          task_stealSide_taskOut_24_TREADY,
  output         task_stealSide_taskOut_24_TVALID,
  output [255:0] task_stealSide_taskOut_24_TDATA,
  input          task_stealSide_taskOut_25_TREADY,
  output         task_stealSide_taskOut_25_TVALID,
  output [255:0] task_stealSide_taskOut_25_TDATA,
  input          task_stealSide_taskOut_26_TREADY,
  output         task_stealSide_taskOut_26_TVALID,
  output [255:0] task_stealSide_taskOut_26_TDATA,
  input          task_stealSide_taskOut_27_TREADY,
  output         task_stealSide_taskOut_27_TVALID,
  output [255:0] task_stealSide_taskOut_27_TDATA,
  input          task_stealSide_taskOut_28_TREADY,
  output         task_stealSide_taskOut_28_TVALID,
  output [255:0] task_stealSide_taskOut_28_TDATA,
  input          task_stealSide_taskOut_29_TREADY,
  output         task_stealSide_taskOut_29_TVALID,
  output [255:0] task_stealSide_taskOut_29_TDATA,
  input          task_stealSide_taskOut_30_TREADY,
  output         task_stealSide_taskOut_30_TVALID,
  output [255:0] task_stealSide_taskOut_30_TDATA,
  input          task_stealSide_taskOut_31_TREADY,
  output         task_stealSide_taskOut_31_TVALID,
  output [255:0] task_stealSide_taskOut_31_TDATA,
  input          task_stealSide_taskOut_32_TREADY,
  output         task_stealSide_taskOut_32_TVALID,
  output [255:0] task_stealSide_taskOut_32_TDATA,
  input          task_stealSide_taskOut_33_TREADY,
  output         task_stealSide_taskOut_33_TVALID,
  output [255:0] task_stealSide_taskOut_33_TDATA,
  input          task_stealSide_taskOut_34_TREADY,
  output         task_stealSide_taskOut_34_TVALID,
  output [255:0] task_stealSide_taskOut_34_TDATA,
  input          task_stealSide_taskOut_35_TREADY,
  output         task_stealSide_taskOut_35_TVALID,
  output [255:0] task_stealSide_taskOut_35_TDATA,
  input          task_stealSide_taskOut_36_TREADY,
  output         task_stealSide_taskOut_36_TVALID,
  output [255:0] task_stealSide_taskOut_36_TDATA,
  input          task_stealSide_taskOut_37_TREADY,
  output         task_stealSide_taskOut_37_TVALID,
  output [255:0] task_stealSide_taskOut_37_TDATA,
  input          task_stealSide_taskOut_38_TREADY,
  output         task_stealSide_taskOut_38_TVALID,
  output [255:0] task_stealSide_taskOut_38_TDATA,
  input          task_stealSide_taskOut_39_TREADY,
  output         task_stealSide_taskOut_39_TVALID,
  output [255:0] task_stealSide_taskOut_39_TDATA,
  input          task_stealSide_taskOut_40_TREADY,
  output         task_stealSide_taskOut_40_TVALID,
  output [255:0] task_stealSide_taskOut_40_TDATA,
  input          task_stealSide_taskOut_41_TREADY,
  output         task_stealSide_taskOut_41_TVALID,
  output [255:0] task_stealSide_taskOut_41_TDATA,
  input          task_stealSide_taskOut_42_TREADY,
  output         task_stealSide_taskOut_42_TVALID,
  output [255:0] task_stealSide_taskOut_42_TDATA,
  input          task_stealSide_taskOut_43_TREADY,
  output         task_stealSide_taskOut_43_TVALID,
  output [255:0] task_stealSide_taskOut_43_TDATA,
  input          task_stealSide_taskOut_44_TREADY,
  output         task_stealSide_taskOut_44_TVALID,
  output [255:0] task_stealSide_taskOut_44_TDATA,
  input          task_stealSide_taskOut_45_TREADY,
  output         task_stealSide_taskOut_45_TVALID,
  output [255:0] task_stealSide_taskOut_45_TDATA,
  input          task_stealSide_taskOut_46_TREADY,
  output         task_stealSide_taskOut_46_TVALID,
  output [255:0] task_stealSide_taskOut_46_TDATA,
  input          task_stealSide_taskOut_47_TREADY,
  output         task_stealSide_taskOut_47_TVALID,
  output [255:0] task_stealSide_taskOut_47_TDATA,
  input          task_stealSide_taskOut_48_TREADY,
  output         task_stealSide_taskOut_48_TVALID,
  output [255:0] task_stealSide_taskOut_48_TDATA,
  input          task_stealSide_taskOut_49_TREADY,
  output         task_stealSide_taskOut_49_TVALID,
  output [255:0] task_stealSide_taskOut_49_TDATA,
  input          task_stealSide_taskOut_50_TREADY,
  output         task_stealSide_taskOut_50_TVALID,
  output [255:0] task_stealSide_taskOut_50_TDATA,
  input          task_stealSide_taskOut_51_TREADY,
  output         task_stealSide_taskOut_51_TVALID,
  output [255:0] task_stealSide_taskOut_51_TDATA,
  input          task_stealSide_taskOut_52_TREADY,
  output         task_stealSide_taskOut_52_TVALID,
  output [255:0] task_stealSide_taskOut_52_TDATA,
  input          task_stealSide_taskOut_53_TREADY,
  output         task_stealSide_taskOut_53_TVALID,
  output [255:0] task_stealSide_taskOut_53_TDATA,
  input          task_stealSide_taskOut_54_TREADY,
  output         task_stealSide_taskOut_54_TVALID,
  output [255:0] task_stealSide_taskOut_54_TDATA,
  input          task_stealSide_taskOut_55_TREADY,
  output         task_stealSide_taskOut_55_TVALID,
  output [255:0] task_stealSide_taskOut_55_TDATA,
  input          task_stealSide_taskOut_56_TREADY,
  output         task_stealSide_taskOut_56_TVALID,
  output [255:0] task_stealSide_taskOut_56_TDATA,
  input          task_stealSide_taskOut_57_TREADY,
  output         task_stealSide_taskOut_57_TVALID,
  output [255:0] task_stealSide_taskOut_57_TDATA,
  input          task_stealSide_taskOut_58_TREADY,
  output         task_stealSide_taskOut_58_TVALID,
  output [255:0] task_stealSide_taskOut_58_TDATA,
  input          task_stealSide_taskOut_59_TREADY,
  output         task_stealSide_taskOut_59_TVALID,
  output [255:0] task_stealSide_taskOut_59_TDATA,
  input          task_stealSide_taskOut_60_TREADY,
  output         task_stealSide_taskOut_60_TVALID,
  output [255:0] task_stealSide_taskOut_60_TDATA,
  input          task_stealSide_taskOut_61_TREADY,
  output         task_stealSide_taskOut_61_TVALID,
  output [255:0] task_stealSide_taskOut_61_TDATA,
  input          task_stealSide_taskOut_62_TREADY,
  output         task_stealSide_taskOut_62_TVALID,
  output [255:0] task_stealSide_taskOut_62_TDATA,
  input          task_stealSide_taskOut_63_TREADY,
  output         task_stealSide_taskOut_63_TVALID,
  output [255:0] task_stealSide_taskOut_63_TDATA,
  output         task_stealSide_taskIn_0_TREADY,
  input          task_stealSide_taskIn_0_TVALID,
  input  [255:0] task_stealSide_taskIn_0_TDATA,
  output         task_stealSide_taskIn_1_TREADY,
  input          task_stealSide_taskIn_1_TVALID,
  input  [255:0] task_stealSide_taskIn_1_TDATA,
  output         task_stealSide_taskIn_2_TREADY,
  input          task_stealSide_taskIn_2_TVALID,
  input  [255:0] task_stealSide_taskIn_2_TDATA,
  output         task_stealSide_taskIn_3_TREADY,
  input          task_stealSide_taskIn_3_TVALID,
  input  [255:0] task_stealSide_taskIn_3_TDATA,
  output         task_stealSide_taskIn_4_TREADY,
  input          task_stealSide_taskIn_4_TVALID,
  input  [255:0] task_stealSide_taskIn_4_TDATA,
  output         task_stealSide_taskIn_5_TREADY,
  input          task_stealSide_taskIn_5_TVALID,
  input  [255:0] task_stealSide_taskIn_5_TDATA,
  output         task_stealSide_taskIn_6_TREADY,
  input          task_stealSide_taskIn_6_TVALID,
  input  [255:0] task_stealSide_taskIn_6_TDATA,
  output         task_stealSide_taskIn_7_TREADY,
  input          task_stealSide_taskIn_7_TVALID,
  input  [255:0] task_stealSide_taskIn_7_TDATA,
  output         task_stealSide_taskIn_8_TREADY,
  input          task_stealSide_taskIn_8_TVALID,
  input  [255:0] task_stealSide_taskIn_8_TDATA,
  output         task_stealSide_taskIn_9_TREADY,
  input          task_stealSide_taskIn_9_TVALID,
  input  [255:0] task_stealSide_taskIn_9_TDATA,
  output         task_stealSide_taskIn_10_TREADY,
  input          task_stealSide_taskIn_10_TVALID,
  input  [255:0] task_stealSide_taskIn_10_TDATA,
  output         task_stealSide_taskIn_11_TREADY,
  input          task_stealSide_taskIn_11_TVALID,
  input  [255:0] task_stealSide_taskIn_11_TDATA,
  output         task_stealSide_taskIn_12_TREADY,
  input          task_stealSide_taskIn_12_TVALID,
  input  [255:0] task_stealSide_taskIn_12_TDATA,
  output         task_stealSide_taskIn_13_TREADY,
  input          task_stealSide_taskIn_13_TVALID,
  input  [255:0] task_stealSide_taskIn_13_TDATA,
  output         task_stealSide_taskIn_14_TREADY,
  input          task_stealSide_taskIn_14_TVALID,
  input  [255:0] task_stealSide_taskIn_14_TDATA,
  output         task_stealSide_taskIn_15_TREADY,
  input          task_stealSide_taskIn_15_TVALID,
  input  [255:0] task_stealSide_taskIn_15_TDATA,
  output         task_stealSide_taskIn_16_TREADY,
  input          task_stealSide_taskIn_16_TVALID,
  input  [255:0] task_stealSide_taskIn_16_TDATA,
  output         task_stealSide_taskIn_17_TREADY,
  input          task_stealSide_taskIn_17_TVALID,
  input  [255:0] task_stealSide_taskIn_17_TDATA,
  output         task_stealSide_taskIn_18_TREADY,
  input          task_stealSide_taskIn_18_TVALID,
  input  [255:0] task_stealSide_taskIn_18_TDATA,
  output         task_stealSide_taskIn_19_TREADY,
  input          task_stealSide_taskIn_19_TVALID,
  input  [255:0] task_stealSide_taskIn_19_TDATA,
  output         task_stealSide_taskIn_20_TREADY,
  input          task_stealSide_taskIn_20_TVALID,
  input  [255:0] task_stealSide_taskIn_20_TDATA,
  output         task_stealSide_taskIn_21_TREADY,
  input          task_stealSide_taskIn_21_TVALID,
  input  [255:0] task_stealSide_taskIn_21_TDATA,
  output         task_stealSide_taskIn_22_TREADY,
  input          task_stealSide_taskIn_22_TVALID,
  input  [255:0] task_stealSide_taskIn_22_TDATA,
  output         task_stealSide_taskIn_23_TREADY,
  input          task_stealSide_taskIn_23_TVALID,
  input  [255:0] task_stealSide_taskIn_23_TDATA,
  output         task_stealSide_taskIn_24_TREADY,
  input          task_stealSide_taskIn_24_TVALID,
  input  [255:0] task_stealSide_taskIn_24_TDATA,
  output         task_stealSide_taskIn_25_TREADY,
  input          task_stealSide_taskIn_25_TVALID,
  input  [255:0] task_stealSide_taskIn_25_TDATA,
  output         task_stealSide_taskIn_26_TREADY,
  input          task_stealSide_taskIn_26_TVALID,
  input  [255:0] task_stealSide_taskIn_26_TDATA,
  output         task_stealSide_taskIn_27_TREADY,
  input          task_stealSide_taskIn_27_TVALID,
  input  [255:0] task_stealSide_taskIn_27_TDATA,
  output         task_stealSide_taskIn_28_TREADY,
  input          task_stealSide_taskIn_28_TVALID,
  input  [255:0] task_stealSide_taskIn_28_TDATA,
  output         task_stealSide_taskIn_29_TREADY,
  input          task_stealSide_taskIn_29_TVALID,
  input  [255:0] task_stealSide_taskIn_29_TDATA,
  output         task_stealSide_taskIn_30_TREADY,
  input          task_stealSide_taskIn_30_TVALID,
  input  [255:0] task_stealSide_taskIn_30_TDATA,
  output         task_stealSide_taskIn_31_TREADY,
  input          task_stealSide_taskIn_31_TVALID,
  input  [255:0] task_stealSide_taskIn_31_TDATA,
  output         task_stealSide_taskIn_32_TREADY,
  input          task_stealSide_taskIn_32_TVALID,
  input  [255:0] task_stealSide_taskIn_32_TDATA,
  output         task_stealSide_taskIn_33_TREADY,
  input          task_stealSide_taskIn_33_TVALID,
  input  [255:0] task_stealSide_taskIn_33_TDATA,
  output         task_stealSide_taskIn_34_TREADY,
  input          task_stealSide_taskIn_34_TVALID,
  input  [255:0] task_stealSide_taskIn_34_TDATA,
  output         task_stealSide_taskIn_35_TREADY,
  input          task_stealSide_taskIn_35_TVALID,
  input  [255:0] task_stealSide_taskIn_35_TDATA,
  output         task_stealSide_taskIn_36_TREADY,
  input          task_stealSide_taskIn_36_TVALID,
  input  [255:0] task_stealSide_taskIn_36_TDATA,
  output         task_stealSide_taskIn_37_TREADY,
  input          task_stealSide_taskIn_37_TVALID,
  input  [255:0] task_stealSide_taskIn_37_TDATA,
  output         task_stealSide_taskIn_38_TREADY,
  input          task_stealSide_taskIn_38_TVALID,
  input  [255:0] task_stealSide_taskIn_38_TDATA,
  output         task_stealSide_taskIn_39_TREADY,
  input          task_stealSide_taskIn_39_TVALID,
  input  [255:0] task_stealSide_taskIn_39_TDATA,
  output         task_stealSide_taskIn_40_TREADY,
  input          task_stealSide_taskIn_40_TVALID,
  input  [255:0] task_stealSide_taskIn_40_TDATA,
  output         task_stealSide_taskIn_41_TREADY,
  input          task_stealSide_taskIn_41_TVALID,
  input  [255:0] task_stealSide_taskIn_41_TDATA,
  output         task_stealSide_taskIn_42_TREADY,
  input          task_stealSide_taskIn_42_TVALID,
  input  [255:0] task_stealSide_taskIn_42_TDATA,
  output         task_stealSide_taskIn_43_TREADY,
  input          task_stealSide_taskIn_43_TVALID,
  input  [255:0] task_stealSide_taskIn_43_TDATA,
  output         task_stealSide_taskIn_44_TREADY,
  input          task_stealSide_taskIn_44_TVALID,
  input  [255:0] task_stealSide_taskIn_44_TDATA,
  output         task_stealSide_taskIn_45_TREADY,
  input          task_stealSide_taskIn_45_TVALID,
  input  [255:0] task_stealSide_taskIn_45_TDATA,
  output         task_stealSide_taskIn_46_TREADY,
  input          task_stealSide_taskIn_46_TVALID,
  input  [255:0] task_stealSide_taskIn_46_TDATA,
  output         task_stealSide_taskIn_47_TREADY,
  input          task_stealSide_taskIn_47_TVALID,
  input  [255:0] task_stealSide_taskIn_47_TDATA,
  output         task_stealSide_taskIn_48_TREADY,
  input          task_stealSide_taskIn_48_TVALID,
  input  [255:0] task_stealSide_taskIn_48_TDATA,
  output         task_stealSide_taskIn_49_TREADY,
  input          task_stealSide_taskIn_49_TVALID,
  input  [255:0] task_stealSide_taskIn_49_TDATA,
  output         task_stealSide_taskIn_50_TREADY,
  input          task_stealSide_taskIn_50_TVALID,
  input  [255:0] task_stealSide_taskIn_50_TDATA,
  output         task_stealSide_taskIn_51_TREADY,
  input          task_stealSide_taskIn_51_TVALID,
  input  [255:0] task_stealSide_taskIn_51_TDATA,
  output         task_stealSide_taskIn_52_TREADY,
  input          task_stealSide_taskIn_52_TVALID,
  input  [255:0] task_stealSide_taskIn_52_TDATA,
  output         task_stealSide_taskIn_53_TREADY,
  input          task_stealSide_taskIn_53_TVALID,
  input  [255:0] task_stealSide_taskIn_53_TDATA,
  output         task_stealSide_taskIn_54_TREADY,
  input          task_stealSide_taskIn_54_TVALID,
  input  [255:0] task_stealSide_taskIn_54_TDATA,
  output         task_stealSide_taskIn_55_TREADY,
  input          task_stealSide_taskIn_55_TVALID,
  input  [255:0] task_stealSide_taskIn_55_TDATA,
  output         task_stealSide_taskIn_56_TREADY,
  input          task_stealSide_taskIn_56_TVALID,
  input  [255:0] task_stealSide_taskIn_56_TDATA,
  output         task_stealSide_taskIn_57_TREADY,
  input          task_stealSide_taskIn_57_TVALID,
  input  [255:0] task_stealSide_taskIn_57_TDATA,
  output         task_stealSide_taskIn_58_TREADY,
  input          task_stealSide_taskIn_58_TVALID,
  input  [255:0] task_stealSide_taskIn_58_TDATA,
  output         task_stealSide_taskIn_59_TREADY,
  input          task_stealSide_taskIn_59_TVALID,
  input  [255:0] task_stealSide_taskIn_59_TDATA,
  output         task_stealSide_taskIn_60_TREADY,
  input          task_stealSide_taskIn_60_TVALID,
  input  [255:0] task_stealSide_taskIn_60_TDATA,
  output         task_stealSide_taskIn_61_TREADY,
  input          task_stealSide_taskIn_61_TVALID,
  input  [255:0] task_stealSide_taskIn_61_TDATA,
  output         task_stealSide_taskIn_62_TREADY,
  input          task_stealSide_taskIn_62_TVALID,
  input  [255:0] task_stealSide_taskIn_62_TDATA,
  output         task_stealSide_taskIn_63_TREADY,
  input          task_stealSide_taskIn_63_TVALID,
  input  [255:0] task_stealSide_taskIn_63_TDATA,
  input          task_continuationAllocationSide_contOut_0_TREADY,
  output         task_continuationAllocationSide_contOut_0_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_0_TDATA,
  input          task_continuationAllocationSide_contOut_1_TREADY,
  output         task_continuationAllocationSide_contOut_1_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_1_TDATA,
  input          task_continuationAllocationSide_contOut_2_TREADY,
  output         task_continuationAllocationSide_contOut_2_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_2_TDATA,
  input          task_continuationAllocationSide_contOut_3_TREADY,
  output         task_continuationAllocationSide_contOut_3_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_3_TDATA,
  input          task_continuationAllocationSide_contOut_4_TREADY,
  output         task_continuationAllocationSide_contOut_4_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_4_TDATA,
  input          task_continuationAllocationSide_contOut_5_TREADY,
  output         task_continuationAllocationSide_contOut_5_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_5_TDATA,
  input          task_continuationAllocationSide_contOut_6_TREADY,
  output         task_continuationAllocationSide_contOut_6_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_6_TDATA,
  input          task_continuationAllocationSide_contOut_7_TREADY,
  output         task_continuationAllocationSide_contOut_7_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_7_TDATA,
  input          task_continuationAllocationSide_contOut_8_TREADY,
  output         task_continuationAllocationSide_contOut_8_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_8_TDATA,
  input          task_continuationAllocationSide_contOut_9_TREADY,
  output         task_continuationAllocationSide_contOut_9_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_9_TDATA,
  input          task_continuationAllocationSide_contOut_10_TREADY,
  output         task_continuationAllocationSide_contOut_10_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_10_TDATA,
  input          task_continuationAllocationSide_contOut_11_TREADY,
  output         task_continuationAllocationSide_contOut_11_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_11_TDATA,
  input          task_continuationAllocationSide_contOut_12_TREADY,
  output         task_continuationAllocationSide_contOut_12_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_12_TDATA,
  input          task_continuationAllocationSide_contOut_13_TREADY,
  output         task_continuationAllocationSide_contOut_13_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_13_TDATA,
  input          task_continuationAllocationSide_contOut_14_TREADY,
  output         task_continuationAllocationSide_contOut_14_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_14_TDATA,
  input          task_continuationAllocationSide_contOut_15_TREADY,
  output         task_continuationAllocationSide_contOut_15_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_15_TDATA,
  input          task_continuationAllocationSide_contOut_16_TREADY,
  output         task_continuationAllocationSide_contOut_16_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_16_TDATA,
  input          task_continuationAllocationSide_contOut_17_TREADY,
  output         task_continuationAllocationSide_contOut_17_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_17_TDATA,
  input          task_continuationAllocationSide_contOut_18_TREADY,
  output         task_continuationAllocationSide_contOut_18_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_18_TDATA,
  input          task_continuationAllocationSide_contOut_19_TREADY,
  output         task_continuationAllocationSide_contOut_19_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_19_TDATA,
  input          task_continuationAllocationSide_contOut_20_TREADY,
  output         task_continuationAllocationSide_contOut_20_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_20_TDATA,
  input          task_continuationAllocationSide_contOut_21_TREADY,
  output         task_continuationAllocationSide_contOut_21_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_21_TDATA,
  input          task_continuationAllocationSide_contOut_22_TREADY,
  output         task_continuationAllocationSide_contOut_22_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_22_TDATA,
  input          task_continuationAllocationSide_contOut_23_TREADY,
  output         task_continuationAllocationSide_contOut_23_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_23_TDATA,
  input          task_continuationAllocationSide_contOut_24_TREADY,
  output         task_continuationAllocationSide_contOut_24_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_24_TDATA,
  input          task_continuationAllocationSide_contOut_25_TREADY,
  output         task_continuationAllocationSide_contOut_25_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_25_TDATA,
  input          task_continuationAllocationSide_contOut_26_TREADY,
  output         task_continuationAllocationSide_contOut_26_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_26_TDATA,
  input          task_continuationAllocationSide_contOut_27_TREADY,
  output         task_continuationAllocationSide_contOut_27_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_27_TDATA,
  input          task_continuationAllocationSide_contOut_28_TREADY,
  output         task_continuationAllocationSide_contOut_28_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_28_TDATA,
  input          task_continuationAllocationSide_contOut_29_TREADY,
  output         task_continuationAllocationSide_contOut_29_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_29_TDATA,
  input          task_continuationAllocationSide_contOut_30_TREADY,
  output         task_continuationAllocationSide_contOut_30_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_30_TDATA,
  input          task_continuationAllocationSide_contOut_31_TREADY,
  output         task_continuationAllocationSide_contOut_31_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_31_TDATA,
  input          task_continuationAllocationSide_contOut_32_TREADY,
  output         task_continuationAllocationSide_contOut_32_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_32_TDATA,
  input          task_continuationAllocationSide_contOut_33_TREADY,
  output         task_continuationAllocationSide_contOut_33_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_33_TDATA,
  input          task_continuationAllocationSide_contOut_34_TREADY,
  output         task_continuationAllocationSide_contOut_34_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_34_TDATA,
  input          task_continuationAllocationSide_contOut_35_TREADY,
  output         task_continuationAllocationSide_contOut_35_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_35_TDATA,
  input          task_continuationAllocationSide_contOut_36_TREADY,
  output         task_continuationAllocationSide_contOut_36_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_36_TDATA,
  input          task_continuationAllocationSide_contOut_37_TREADY,
  output         task_continuationAllocationSide_contOut_37_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_37_TDATA,
  input          task_continuationAllocationSide_contOut_38_TREADY,
  output         task_continuationAllocationSide_contOut_38_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_38_TDATA,
  input          task_continuationAllocationSide_contOut_39_TREADY,
  output         task_continuationAllocationSide_contOut_39_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_39_TDATA,
  input          task_continuationAllocationSide_contOut_40_TREADY,
  output         task_continuationAllocationSide_contOut_40_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_40_TDATA,
  input          task_continuationAllocationSide_contOut_41_TREADY,
  output         task_continuationAllocationSide_contOut_41_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_41_TDATA,
  input          task_continuationAllocationSide_contOut_42_TREADY,
  output         task_continuationAllocationSide_contOut_42_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_42_TDATA,
  input          task_continuationAllocationSide_contOut_43_TREADY,
  output         task_continuationAllocationSide_contOut_43_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_43_TDATA,
  input          task_continuationAllocationSide_contOut_44_TREADY,
  output         task_continuationAllocationSide_contOut_44_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_44_TDATA,
  input          task_continuationAllocationSide_contOut_45_TREADY,
  output         task_continuationAllocationSide_contOut_45_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_45_TDATA,
  input          task_continuationAllocationSide_contOut_46_TREADY,
  output         task_continuationAllocationSide_contOut_46_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_46_TDATA,
  input          task_continuationAllocationSide_contOut_47_TREADY,
  output         task_continuationAllocationSide_contOut_47_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_47_TDATA,
  input          task_continuationAllocationSide_contOut_48_TREADY,
  output         task_continuationAllocationSide_contOut_48_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_48_TDATA,
  input          task_continuationAllocationSide_contOut_49_TREADY,
  output         task_continuationAllocationSide_contOut_49_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_49_TDATA,
  input          task_continuationAllocationSide_contOut_50_TREADY,
  output         task_continuationAllocationSide_contOut_50_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_50_TDATA,
  input          task_continuationAllocationSide_contOut_51_TREADY,
  output         task_continuationAllocationSide_contOut_51_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_51_TDATA,
  input          task_continuationAllocationSide_contOut_52_TREADY,
  output         task_continuationAllocationSide_contOut_52_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_52_TDATA,
  input          task_continuationAllocationSide_contOut_53_TREADY,
  output         task_continuationAllocationSide_contOut_53_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_53_TDATA,
  input          task_continuationAllocationSide_contOut_54_TREADY,
  output         task_continuationAllocationSide_contOut_54_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_54_TDATA,
  input          task_continuationAllocationSide_contOut_55_TREADY,
  output         task_continuationAllocationSide_contOut_55_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_55_TDATA,
  input          task_continuationAllocationSide_contOut_56_TREADY,
  output         task_continuationAllocationSide_contOut_56_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_56_TDATA,
  input          task_continuationAllocationSide_contOut_57_TREADY,
  output         task_continuationAllocationSide_contOut_57_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_57_TDATA,
  input          task_continuationAllocationSide_contOut_58_TREADY,
  output         task_continuationAllocationSide_contOut_58_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_58_TDATA,
  input          task_continuationAllocationSide_contOut_59_TREADY,
  output         task_continuationAllocationSide_contOut_59_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_59_TDATA,
  input          task_continuationAllocationSide_contOut_60_TREADY,
  output         task_continuationAllocationSide_contOut_60_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_60_TDATA,
  input          task_continuationAllocationSide_contOut_61_TREADY,
  output         task_continuationAllocationSide_contOut_61_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_61_TDATA,
  input          task_continuationAllocationSide_contOut_62_TREADY,
  output         task_continuationAllocationSide_contOut_62_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_62_TDATA,
  input          task_continuationAllocationSide_contOut_63_TREADY,
  output         task_continuationAllocationSide_contOut_63_TVALID,
  output [63:0]  task_continuationAllocationSide_contOut_63_TDATA,
  output         task_continuationAllocationSide_axi_mgmt_vcas_0_ARREADY,
  input          task_continuationAllocationSide_axi_mgmt_vcas_0_ARVALID,
  input  [5:0]   task_continuationAllocationSide_axi_mgmt_vcas_0_ARADDR,
  input  [2:0]   task_continuationAllocationSide_axi_mgmt_vcas_0_ARPROT,
  input          task_continuationAllocationSide_axi_mgmt_vcas_0_RREADY,
  output         task_continuationAllocationSide_axi_mgmt_vcas_0_RVALID,
  output [63:0]  task_continuationAllocationSide_axi_mgmt_vcas_0_RDATA,
  output [1:0]   task_continuationAllocationSide_axi_mgmt_vcas_0_RRESP,
  output         task_continuationAllocationSide_axi_mgmt_vcas_0_AWREADY,
  input          task_continuationAllocationSide_axi_mgmt_vcas_0_AWVALID,
  input  [5:0]   task_continuationAllocationSide_axi_mgmt_vcas_0_AWADDR,
  input  [2:0]   task_continuationAllocationSide_axi_mgmt_vcas_0_AWPROT,
  output         task_continuationAllocationSide_axi_mgmt_vcas_0_WREADY,
  input          task_continuationAllocationSide_axi_mgmt_vcas_0_WVALID,
  input  [63:0]  task_continuationAllocationSide_axi_mgmt_vcas_0_WDATA,
  input  [7:0]   task_continuationAllocationSide_axi_mgmt_vcas_0_WSTRB,
  input          task_continuationAllocationSide_axi_mgmt_vcas_0_BREADY,
  output         task_continuationAllocationSide_axi_mgmt_vcas_0_BVALID,
  output [1:0]   task_continuationAllocationSide_axi_mgmt_vcas_0_BRESP,
  input          task_continuationAllocationSide_vcas_axi_full_0_ARREADY,
  output         task_continuationAllocationSide_vcas_axi_full_0_ARVALID,
  output [3:0]   task_continuationAllocationSide_vcas_axi_full_0_ARID,
  output [63:0]  task_continuationAllocationSide_vcas_axi_full_0_ARADDR,
  output [7:0]   task_continuationAllocationSide_vcas_axi_full_0_ARLEN,
  output [2:0]   task_continuationAllocationSide_vcas_axi_full_0_ARSIZE,
  output [1:0]   task_continuationAllocationSide_vcas_axi_full_0_ARBURST,
  output         task_continuationAllocationSide_vcas_axi_full_0_ARLOCK,
  output [3:0]   task_continuationAllocationSide_vcas_axi_full_0_ARCACHE,
  output [2:0]   task_continuationAllocationSide_vcas_axi_full_0_ARPROT,
  output [3:0]   task_continuationAllocationSide_vcas_axi_full_0_ARQOS,
  output [3:0]   task_continuationAllocationSide_vcas_axi_full_0_ARREGION,
  output         task_continuationAllocationSide_vcas_axi_full_0_RREADY,
  input          task_continuationAllocationSide_vcas_axi_full_0_RVALID,
  input  [3:0]   task_continuationAllocationSide_vcas_axi_full_0_RID,
  input  [63:0]  task_continuationAllocationSide_vcas_axi_full_0_RDATA,
  input  [1:0]   task_continuationAllocationSide_vcas_axi_full_0_RRESP,
  input          task_continuationAllocationSide_vcas_axi_full_0_RLAST,
  input          task_continuationAllocationSide_vcas_axi_full_0_AWREADY,
  output         task_continuationAllocationSide_vcas_axi_full_0_AWVALID,
  output [3:0]   task_continuationAllocationSide_vcas_axi_full_0_AWID,
  output [63:0]  task_continuationAllocationSide_vcas_axi_full_0_AWADDR,
  output [7:0]   task_continuationAllocationSide_vcas_axi_full_0_AWLEN,
  output [2:0]   task_continuationAllocationSide_vcas_axi_full_0_AWSIZE,
  output [1:0]   task_continuationAllocationSide_vcas_axi_full_0_AWBURST,
  output         task_continuationAllocationSide_vcas_axi_full_0_AWLOCK,
  output [3:0]   task_continuationAllocationSide_vcas_axi_full_0_AWCACHE,
  output [2:0]   task_continuationAllocationSide_vcas_axi_full_0_AWPROT,
  output [3:0]   task_continuationAllocationSide_vcas_axi_full_0_AWQOS,
  output [3:0]   task_continuationAllocationSide_vcas_axi_full_0_AWREGION,
  input          task_continuationAllocationSide_vcas_axi_full_0_WREADY,
  output         task_continuationAllocationSide_vcas_axi_full_0_WVALID,
  output [3:0]   task_continuationAllocationSide_vcas_axi_full_0_WID,
  output [63:0]  task_continuationAllocationSide_vcas_axi_full_0_WDATA,
  output [7:0]   task_continuationAllocationSide_vcas_axi_full_0_WSTRB,
  output         task_continuationAllocationSide_vcas_axi_full_0_WLAST,
  output         task_continuationAllocationSide_vcas_axi_full_0_BREADY,
  input          task_continuationAllocationSide_vcas_axi_full_0_BVALID,
  input  [3:0]   task_continuationAllocationSide_vcas_axi_full_0_BID,
  input  [1:0]   task_continuationAllocationSide_vcas_axi_full_0_BRESP,
  output         task_syncSide_addrIn_0_TREADY,
  input          task_syncSide_addrIn_0_TVALID,
  input  [63:0]  task_syncSide_addrIn_0_TDATA,
  output         task_syncSide_addrIn_1_TREADY,
  input          task_syncSide_addrIn_1_TVALID,
  input  [63:0]  task_syncSide_addrIn_1_TDATA,
  output         task_syncSide_addrIn_2_TREADY,
  input          task_syncSide_addrIn_2_TVALID,
  input  [63:0]  task_syncSide_addrIn_2_TDATA,
  output         task_syncSide_addrIn_3_TREADY,
  input          task_syncSide_addrIn_3_TVALID,
  input  [63:0]  task_syncSide_addrIn_3_TDATA,
  output         task_syncSide_addrIn_4_TREADY,
  input          task_syncSide_addrIn_4_TVALID,
  input  [63:0]  task_syncSide_addrIn_4_TDATA,
  output         task_syncSide_addrIn_5_TREADY,
  input          task_syncSide_addrIn_5_TVALID,
  input  [63:0]  task_syncSide_addrIn_5_TDATA,
  output         task_syncSide_addrIn_6_TREADY,
  input          task_syncSide_addrIn_6_TVALID,
  input  [63:0]  task_syncSide_addrIn_6_TDATA,
  output         task_syncSide_addrIn_7_TREADY,
  input          task_syncSide_addrIn_7_TVALID,
  input  [63:0]  task_syncSide_addrIn_7_TDATA,
  output         task_syncSide_addrIn_8_TREADY,
  input          task_syncSide_addrIn_8_TVALID,
  input  [63:0]  task_syncSide_addrIn_8_TDATA,
  output         task_syncSide_addrIn_9_TREADY,
  input          task_syncSide_addrIn_9_TVALID,
  input  [63:0]  task_syncSide_addrIn_9_TDATA,
  output         task_syncSide_addrIn_10_TREADY,
  input          task_syncSide_addrIn_10_TVALID,
  input  [63:0]  task_syncSide_addrIn_10_TDATA,
  output         task_syncSide_addrIn_11_TREADY,
  input          task_syncSide_addrIn_11_TVALID,
  input  [63:0]  task_syncSide_addrIn_11_TDATA,
  output         task_syncSide_addrIn_12_TREADY,
  input          task_syncSide_addrIn_12_TVALID,
  input  [63:0]  task_syncSide_addrIn_12_TDATA,
  output         task_syncSide_addrIn_13_TREADY,
  input          task_syncSide_addrIn_13_TVALID,
  input  [63:0]  task_syncSide_addrIn_13_TDATA,
  output         task_syncSide_addrIn_14_TREADY,
  input          task_syncSide_addrIn_14_TVALID,
  input  [63:0]  task_syncSide_addrIn_14_TDATA,
  output         task_syncSide_addrIn_15_TREADY,
  input          task_syncSide_addrIn_15_TVALID,
  input  [63:0]  task_syncSide_addrIn_15_TDATA,
  output         task_syncSide_addrIn_16_TREADY,
  input          task_syncSide_addrIn_16_TVALID,
  input  [63:0]  task_syncSide_addrIn_16_TDATA,
  output         task_syncSide_addrIn_17_TREADY,
  input          task_syncSide_addrIn_17_TVALID,
  input  [63:0]  task_syncSide_addrIn_17_TDATA,
  output         task_syncSide_addrIn_18_TREADY,
  input          task_syncSide_addrIn_18_TVALID,
  input  [63:0]  task_syncSide_addrIn_18_TDATA,
  output         task_syncSide_addrIn_19_TREADY,
  input          task_syncSide_addrIn_19_TVALID,
  input  [63:0]  task_syncSide_addrIn_19_TDATA,
  output         task_syncSide_addrIn_20_TREADY,
  input          task_syncSide_addrIn_20_TVALID,
  input  [63:0]  task_syncSide_addrIn_20_TDATA,
  output         task_syncSide_addrIn_21_TREADY,
  input          task_syncSide_addrIn_21_TVALID,
  input  [63:0]  task_syncSide_addrIn_21_TDATA,
  output         task_syncSide_addrIn_22_TREADY,
  input          task_syncSide_addrIn_22_TVALID,
  input  [63:0]  task_syncSide_addrIn_22_TDATA,
  output         task_syncSide_addrIn_23_TREADY,
  input          task_syncSide_addrIn_23_TVALID,
  input  [63:0]  task_syncSide_addrIn_23_TDATA,
  output         task_syncSide_addrIn_24_TREADY,
  input          task_syncSide_addrIn_24_TVALID,
  input  [63:0]  task_syncSide_addrIn_24_TDATA,
  output         task_syncSide_addrIn_25_TREADY,
  input          task_syncSide_addrIn_25_TVALID,
  input  [63:0]  task_syncSide_addrIn_25_TDATA,
  output         task_syncSide_addrIn_26_TREADY,
  input          task_syncSide_addrIn_26_TVALID,
  input  [63:0]  task_syncSide_addrIn_26_TDATA,
  output         task_syncSide_addrIn_27_TREADY,
  input          task_syncSide_addrIn_27_TVALID,
  input  [63:0]  task_syncSide_addrIn_27_TDATA,
  output         task_syncSide_addrIn_28_TREADY,
  input          task_syncSide_addrIn_28_TVALID,
  input  [63:0]  task_syncSide_addrIn_28_TDATA,
  output         task_syncSide_addrIn_29_TREADY,
  input          task_syncSide_addrIn_29_TVALID,
  input  [63:0]  task_syncSide_addrIn_29_TDATA,
  output         task_syncSide_addrIn_30_TREADY,
  input          task_syncSide_addrIn_30_TVALID,
  input  [63:0]  task_syncSide_addrIn_30_TDATA,
  output         task_syncSide_addrIn_31_TREADY,
  input          task_syncSide_addrIn_31_TVALID,
  input  [63:0]  task_syncSide_addrIn_31_TDATA,
  output         task_syncSide_addrIn_32_TREADY,
  input          task_syncSide_addrIn_32_TVALID,
  input  [63:0]  task_syncSide_addrIn_32_TDATA,
  output         task_syncSide_addrIn_33_TREADY,
  input          task_syncSide_addrIn_33_TVALID,
  input  [63:0]  task_syncSide_addrIn_33_TDATA,
  output         task_syncSide_addrIn_34_TREADY,
  input          task_syncSide_addrIn_34_TVALID,
  input  [63:0]  task_syncSide_addrIn_34_TDATA,
  output         task_syncSide_addrIn_35_TREADY,
  input          task_syncSide_addrIn_35_TVALID,
  input  [63:0]  task_syncSide_addrIn_35_TDATA,
  output         task_syncSide_addrIn_36_TREADY,
  input          task_syncSide_addrIn_36_TVALID,
  input  [63:0]  task_syncSide_addrIn_36_TDATA,
  output         task_syncSide_addrIn_37_TREADY,
  input          task_syncSide_addrIn_37_TVALID,
  input  [63:0]  task_syncSide_addrIn_37_TDATA,
  output         task_syncSide_addrIn_38_TREADY,
  input          task_syncSide_addrIn_38_TVALID,
  input  [63:0]  task_syncSide_addrIn_38_TDATA,
  output         task_syncSide_addrIn_39_TREADY,
  input          task_syncSide_addrIn_39_TVALID,
  input  [63:0]  task_syncSide_addrIn_39_TDATA,
  output         task_syncSide_addrIn_40_TREADY,
  input          task_syncSide_addrIn_40_TVALID,
  input  [63:0]  task_syncSide_addrIn_40_TDATA,
  output         task_syncSide_addrIn_41_TREADY,
  input          task_syncSide_addrIn_41_TVALID,
  input  [63:0]  task_syncSide_addrIn_41_TDATA,
  output         task_syncSide_addrIn_42_TREADY,
  input          task_syncSide_addrIn_42_TVALID,
  input  [63:0]  task_syncSide_addrIn_42_TDATA,
  output         task_syncSide_addrIn_43_TREADY,
  input          task_syncSide_addrIn_43_TVALID,
  input  [63:0]  task_syncSide_addrIn_43_TDATA,
  output         task_syncSide_addrIn_44_TREADY,
  input          task_syncSide_addrIn_44_TVALID,
  input  [63:0]  task_syncSide_addrIn_44_TDATA,
  output         task_syncSide_addrIn_45_TREADY,
  input          task_syncSide_addrIn_45_TVALID,
  input  [63:0]  task_syncSide_addrIn_45_TDATA,
  output         task_syncSide_addrIn_46_TREADY,
  input          task_syncSide_addrIn_46_TVALID,
  input  [63:0]  task_syncSide_addrIn_46_TDATA,
  output         task_syncSide_addrIn_47_TREADY,
  input          task_syncSide_addrIn_47_TVALID,
  input  [63:0]  task_syncSide_addrIn_47_TDATA,
  output         task_syncSide_addrIn_48_TREADY,
  input          task_syncSide_addrIn_48_TVALID,
  input  [63:0]  task_syncSide_addrIn_48_TDATA,
  output         task_syncSide_addrIn_49_TREADY,
  input          task_syncSide_addrIn_49_TVALID,
  input  [63:0]  task_syncSide_addrIn_49_TDATA,
  output         task_syncSide_addrIn_50_TREADY,
  input          task_syncSide_addrIn_50_TVALID,
  input  [63:0]  task_syncSide_addrIn_50_TDATA,
  output         task_syncSide_addrIn_51_TREADY,
  input          task_syncSide_addrIn_51_TVALID,
  input  [63:0]  task_syncSide_addrIn_51_TDATA,
  output         task_syncSide_addrIn_52_TREADY,
  input          task_syncSide_addrIn_52_TVALID,
  input  [63:0]  task_syncSide_addrIn_52_TDATA,
  output         task_syncSide_addrIn_53_TREADY,
  input          task_syncSide_addrIn_53_TVALID,
  input  [63:0]  task_syncSide_addrIn_53_TDATA,
  output         task_syncSide_addrIn_54_TREADY,
  input          task_syncSide_addrIn_54_TVALID,
  input  [63:0]  task_syncSide_addrIn_54_TDATA,
  output         task_syncSide_addrIn_55_TREADY,
  input          task_syncSide_addrIn_55_TVALID,
  input  [63:0]  task_syncSide_addrIn_55_TDATA,
  output         task_syncSide_addrIn_56_TREADY,
  input          task_syncSide_addrIn_56_TVALID,
  input  [63:0]  task_syncSide_addrIn_56_TDATA,
  output         task_syncSide_addrIn_57_TREADY,
  input          task_syncSide_addrIn_57_TVALID,
  input  [63:0]  task_syncSide_addrIn_57_TDATA,
  output         task_syncSide_addrIn_58_TREADY,
  input          task_syncSide_addrIn_58_TVALID,
  input  [63:0]  task_syncSide_addrIn_58_TDATA,
  output         task_syncSide_addrIn_59_TREADY,
  input          task_syncSide_addrIn_59_TVALID,
  input  [63:0]  task_syncSide_addrIn_59_TDATA,
  output         task_syncSide_addrIn_60_TREADY,
  input          task_syncSide_addrIn_60_TVALID,
  input  [63:0]  task_syncSide_addrIn_60_TDATA,
  output         task_syncSide_addrIn_61_TREADY,
  input          task_syncSide_addrIn_61_TVALID,
  input  [63:0]  task_syncSide_addrIn_61_TDATA,
  output         task_syncSide_addrIn_62_TREADY,
  input          task_syncSide_addrIn_62_TVALID,
  input  [63:0]  task_syncSide_addrIn_62_TDATA,
  output         task_syncSide_addrIn_63_TREADY,
  input          task_syncSide_addrIn_63_TVALID,
  input  [63:0]  task_syncSide_addrIn_63_TDATA,
  input          task_syncSide_axi_full_argRoute_0_ARREADY,
  output         task_syncSide_axi_full_argRoute_0_ARVALID,
  output [3:0]   task_syncSide_axi_full_argRoute_0_ARID,
  output [63:0]  task_syncSide_axi_full_argRoute_0_ARADDR,
  output [7:0]   task_syncSide_axi_full_argRoute_0_ARLEN,
  output [2:0]   task_syncSide_axi_full_argRoute_0_ARSIZE,
  output [1:0]   task_syncSide_axi_full_argRoute_0_ARBURST,
  output         task_syncSide_axi_full_argRoute_0_ARLOCK,
  output [3:0]   task_syncSide_axi_full_argRoute_0_ARCACHE,
  output [2:0]   task_syncSide_axi_full_argRoute_0_ARPROT,
  output [3:0]   task_syncSide_axi_full_argRoute_0_ARQOS,
  output [3:0]   task_syncSide_axi_full_argRoute_0_ARREGION,
  output         task_syncSide_axi_full_argRoute_0_RREADY,
  input          task_syncSide_axi_full_argRoute_0_RVALID,
  input  [3:0]   task_syncSide_axi_full_argRoute_0_RID,
  input  [31:0]  task_syncSide_axi_full_argRoute_0_RDATA,
  input  [1:0]   task_syncSide_axi_full_argRoute_0_RRESP,
  input          task_syncSide_axi_full_argRoute_0_RLAST,
  input          task_syncSide_axi_full_argRoute_0_AWREADY,
  output         task_syncSide_axi_full_argRoute_0_AWVALID,
  output [3:0]   task_syncSide_axi_full_argRoute_0_AWID,
  output [63:0]  task_syncSide_axi_full_argRoute_0_AWADDR,
  output [7:0]   task_syncSide_axi_full_argRoute_0_AWLEN,
  output [2:0]   task_syncSide_axi_full_argRoute_0_AWSIZE,
  output [1:0]   task_syncSide_axi_full_argRoute_0_AWBURST,
  output         task_syncSide_axi_full_argRoute_0_AWLOCK,
  output [3:0]   task_syncSide_axi_full_argRoute_0_AWCACHE,
  output [2:0]   task_syncSide_axi_full_argRoute_0_AWPROT,
  output [3:0]   task_syncSide_axi_full_argRoute_0_AWQOS,
  output [3:0]   task_syncSide_axi_full_argRoute_0_AWREGION,
  input          task_syncSide_axi_full_argRoute_0_WREADY,
  output         task_syncSide_axi_full_argRoute_0_WVALID,
  output [3:0]   task_syncSide_axi_full_argRoute_0_WID,
  output [31:0]  task_syncSide_axi_full_argRoute_0_WDATA,
  output [3:0]   task_syncSide_axi_full_argRoute_0_WSTRB,
  output         task_syncSide_axi_full_argRoute_0_WLAST,
  output         task_syncSide_axi_full_argRoute_0_BREADY,
  input          task_syncSide_axi_full_argRoute_0_BVALID,
  input  [3:0]   task_syncSide_axi_full_argRoute_0_BID,
  input  [1:0]   task_syncSide_axi_full_argRoute_0_BRESP,
  input          task_syncSide_axi_full_argRoute_1_ARREADY,
  output         task_syncSide_axi_full_argRoute_1_ARVALID,
  output [3:0]   task_syncSide_axi_full_argRoute_1_ARID,
  output [63:0]  task_syncSide_axi_full_argRoute_1_ARADDR,
  output [7:0]   task_syncSide_axi_full_argRoute_1_ARLEN,
  output [2:0]   task_syncSide_axi_full_argRoute_1_ARSIZE,
  output [1:0]   task_syncSide_axi_full_argRoute_1_ARBURST,
  output         task_syncSide_axi_full_argRoute_1_ARLOCK,
  output [3:0]   task_syncSide_axi_full_argRoute_1_ARCACHE,
  output [2:0]   task_syncSide_axi_full_argRoute_1_ARPROT,
  output [3:0]   task_syncSide_axi_full_argRoute_1_ARQOS,
  output [3:0]   task_syncSide_axi_full_argRoute_1_ARREGION,
  output         task_syncSide_axi_full_argRoute_1_RREADY,
  input          task_syncSide_axi_full_argRoute_1_RVALID,
  input  [3:0]   task_syncSide_axi_full_argRoute_1_RID,
  input  [31:0]  task_syncSide_axi_full_argRoute_1_RDATA,
  input  [1:0]   task_syncSide_axi_full_argRoute_1_RRESP,
  input          task_syncSide_axi_full_argRoute_1_RLAST,
  input          task_syncSide_axi_full_argRoute_1_AWREADY,
  output         task_syncSide_axi_full_argRoute_1_AWVALID,
  output [3:0]   task_syncSide_axi_full_argRoute_1_AWID,
  output [63:0]  task_syncSide_axi_full_argRoute_1_AWADDR,
  output [7:0]   task_syncSide_axi_full_argRoute_1_AWLEN,
  output [2:0]   task_syncSide_axi_full_argRoute_1_AWSIZE,
  output [1:0]   task_syncSide_axi_full_argRoute_1_AWBURST,
  output         task_syncSide_axi_full_argRoute_1_AWLOCK,
  output [3:0]   task_syncSide_axi_full_argRoute_1_AWCACHE,
  output [2:0]   task_syncSide_axi_full_argRoute_1_AWPROT,
  output [3:0]   task_syncSide_axi_full_argRoute_1_AWQOS,
  output [3:0]   task_syncSide_axi_full_argRoute_1_AWREGION,
  input          task_syncSide_axi_full_argRoute_1_WREADY,
  output         task_syncSide_axi_full_argRoute_1_WVALID,
  output [3:0]   task_syncSide_axi_full_argRoute_1_WID,
  output [31:0]  task_syncSide_axi_full_argRoute_1_WDATA,
  output [3:0]   task_syncSide_axi_full_argRoute_1_WSTRB,
  output         task_syncSide_axi_full_argRoute_1_WLAST,
  output         task_syncSide_axi_full_argRoute_1_BREADY,
  input          task_syncSide_axi_full_argRoute_1_BVALID,
  input  [3:0]   task_syncSide_axi_full_argRoute_1_BID,
  input  [1:0]   task_syncSide_axi_full_argRoute_1_BRESP,
  input          task_syncSide_axi_full_argRoute_2_ARREADY,
  output         task_syncSide_axi_full_argRoute_2_ARVALID,
  output [3:0]   task_syncSide_axi_full_argRoute_2_ARID,
  output [63:0]  task_syncSide_axi_full_argRoute_2_ARADDR,
  output [7:0]   task_syncSide_axi_full_argRoute_2_ARLEN,
  output [2:0]   task_syncSide_axi_full_argRoute_2_ARSIZE,
  output [1:0]   task_syncSide_axi_full_argRoute_2_ARBURST,
  output         task_syncSide_axi_full_argRoute_2_ARLOCK,
  output [3:0]   task_syncSide_axi_full_argRoute_2_ARCACHE,
  output [2:0]   task_syncSide_axi_full_argRoute_2_ARPROT,
  output [3:0]   task_syncSide_axi_full_argRoute_2_ARQOS,
  output [3:0]   task_syncSide_axi_full_argRoute_2_ARREGION,
  output         task_syncSide_axi_full_argRoute_2_RREADY,
  input          task_syncSide_axi_full_argRoute_2_RVALID,
  input  [3:0]   task_syncSide_axi_full_argRoute_2_RID,
  input  [31:0]  task_syncSide_axi_full_argRoute_2_RDATA,
  input  [1:0]   task_syncSide_axi_full_argRoute_2_RRESP,
  input          task_syncSide_axi_full_argRoute_2_RLAST,
  input          task_syncSide_axi_full_argRoute_2_AWREADY,
  output         task_syncSide_axi_full_argRoute_2_AWVALID,
  output [3:0]   task_syncSide_axi_full_argRoute_2_AWID,
  output [63:0]  task_syncSide_axi_full_argRoute_2_AWADDR,
  output [7:0]   task_syncSide_axi_full_argRoute_2_AWLEN,
  output [2:0]   task_syncSide_axi_full_argRoute_2_AWSIZE,
  output [1:0]   task_syncSide_axi_full_argRoute_2_AWBURST,
  output         task_syncSide_axi_full_argRoute_2_AWLOCK,
  output [3:0]   task_syncSide_axi_full_argRoute_2_AWCACHE,
  output [2:0]   task_syncSide_axi_full_argRoute_2_AWPROT,
  output [3:0]   task_syncSide_axi_full_argRoute_2_AWQOS,
  output [3:0]   task_syncSide_axi_full_argRoute_2_AWREGION,
  input          task_syncSide_axi_full_argRoute_2_WREADY,
  output         task_syncSide_axi_full_argRoute_2_WVALID,
  output [3:0]   task_syncSide_axi_full_argRoute_2_WID,
  output [31:0]  task_syncSide_axi_full_argRoute_2_WDATA,
  output [3:0]   task_syncSide_axi_full_argRoute_2_WSTRB,
  output         task_syncSide_axi_full_argRoute_2_WLAST,
  output         task_syncSide_axi_full_argRoute_2_BREADY,
  input          task_syncSide_axi_full_argRoute_2_BVALID,
  input  [3:0]   task_syncSide_axi_full_argRoute_2_BID,
  input  [1:0]   task_syncSide_axi_full_argRoute_2_BRESP,
  input          task_syncSide_axi_full_argRoute_3_ARREADY,
  output         task_syncSide_axi_full_argRoute_3_ARVALID,
  output [3:0]   task_syncSide_axi_full_argRoute_3_ARID,
  output [63:0]  task_syncSide_axi_full_argRoute_3_ARADDR,
  output [7:0]   task_syncSide_axi_full_argRoute_3_ARLEN,
  output [2:0]   task_syncSide_axi_full_argRoute_3_ARSIZE,
  output [1:0]   task_syncSide_axi_full_argRoute_3_ARBURST,
  output         task_syncSide_axi_full_argRoute_3_ARLOCK,
  output [3:0]   task_syncSide_axi_full_argRoute_3_ARCACHE,
  output [2:0]   task_syncSide_axi_full_argRoute_3_ARPROT,
  output [3:0]   task_syncSide_axi_full_argRoute_3_ARQOS,
  output [3:0]   task_syncSide_axi_full_argRoute_3_ARREGION,
  output         task_syncSide_axi_full_argRoute_3_RREADY,
  input          task_syncSide_axi_full_argRoute_3_RVALID,
  input  [3:0]   task_syncSide_axi_full_argRoute_3_RID,
  input  [31:0]  task_syncSide_axi_full_argRoute_3_RDATA,
  input  [1:0]   task_syncSide_axi_full_argRoute_3_RRESP,
  input          task_syncSide_axi_full_argRoute_3_RLAST,
  input          task_syncSide_axi_full_argRoute_3_AWREADY,
  output         task_syncSide_axi_full_argRoute_3_AWVALID,
  output [3:0]   task_syncSide_axi_full_argRoute_3_AWID,
  output [63:0]  task_syncSide_axi_full_argRoute_3_AWADDR,
  output [7:0]   task_syncSide_axi_full_argRoute_3_AWLEN,
  output [2:0]   task_syncSide_axi_full_argRoute_3_AWSIZE,
  output [1:0]   task_syncSide_axi_full_argRoute_3_AWBURST,
  output         task_syncSide_axi_full_argRoute_3_AWLOCK,
  output [3:0]   task_syncSide_axi_full_argRoute_3_AWCACHE,
  output [2:0]   task_syncSide_axi_full_argRoute_3_AWPROT,
  output [3:0]   task_syncSide_axi_full_argRoute_3_AWQOS,
  output [3:0]   task_syncSide_axi_full_argRoute_3_AWREGION,
  input          task_syncSide_axi_full_argRoute_3_WREADY,
  output         task_syncSide_axi_full_argRoute_3_WVALID,
  output [3:0]   task_syncSide_axi_full_argRoute_3_WID,
  output [31:0]  task_syncSide_axi_full_argRoute_3_WDATA,
  output [3:0]   task_syncSide_axi_full_argRoute_3_WSTRB,
  output         task_syncSide_axi_full_argRoute_3_WLAST,
  output         task_syncSide_axi_full_argRoute_3_BREADY,
  input          task_syncSide_axi_full_argRoute_3_BVALID,
  input  [3:0]   task_syncSide_axi_full_argRoute_3_BID,
  input  [1:0]   task_syncSide_axi_full_argRoute_3_BRESP
);
  wire  stealSide_clock; // @[fullSysGen.scala 228:29]
  wire  stealSide_reset; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_axi_mgmt_vss_0_ARREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_axi_mgmt_vss_0_ARVALID; // @[fullSysGen.scala 228:29]
  wire [5:0] stealSide_io_axi_mgmt_vss_0_ARADDR; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_axi_mgmt_vss_0_RREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_axi_mgmt_vss_0_RVALID; // @[fullSysGen.scala 228:29]
  wire [63:0] stealSide_io_axi_mgmt_vss_0_RDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_axi_mgmt_vss_0_AWREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_axi_mgmt_vss_0_AWVALID; // @[fullSysGen.scala 228:29]
  wire [5:0] stealSide_io_axi_mgmt_vss_0_AWADDR; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_axi_mgmt_vss_0_WREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_axi_mgmt_vss_0_WVALID; // @[fullSysGen.scala 228:29]
  wire [63:0] stealSide_io_axi_mgmt_vss_0_WDATA; // @[fullSysGen.scala 228:29]
  wire [7:0] stealSide_io_axi_mgmt_vss_0_WSTRB; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_axi_mgmt_vss_0_BREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_axi_mgmt_vss_0_BVALID; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_vss_axi_full_0_ARREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_vss_axi_full_0_ARVALID; // @[fullSysGen.scala 228:29]
  wire [63:0] stealSide_io_vss_axi_full_0_ARADDR; // @[fullSysGen.scala 228:29]
  wire [7:0] stealSide_io_vss_axi_full_0_ARLEN; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_vss_axi_full_0_RREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_vss_axi_full_0_RVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_vss_axi_full_0_RDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_vss_axi_full_0_AWREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_vss_axi_full_0_AWVALID; // @[fullSysGen.scala 228:29]
  wire [63:0] stealSide_io_vss_axi_full_0_AWADDR; // @[fullSysGen.scala 228:29]
  wire [7:0] stealSide_io_vss_axi_full_0_AWLEN; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_vss_axi_full_0_WREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_vss_axi_full_0_WVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_vss_axi_full_0_WDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_vss_axi_full_0_WLAST; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_vss_axi_full_0_BVALID; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_0_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_0_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_0_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_1_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_1_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_1_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_2_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_2_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_2_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_3_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_3_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_3_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_4_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_4_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_4_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_5_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_5_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_5_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_6_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_6_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_6_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_7_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_7_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_7_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_8_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_8_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_8_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_9_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_9_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_9_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_10_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_10_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_10_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_11_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_11_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_11_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_12_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_12_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_12_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_13_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_13_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_13_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_14_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_14_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_14_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_15_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_15_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_15_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_16_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_16_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_16_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_17_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_17_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_17_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_18_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_18_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_18_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_19_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_19_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_19_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_20_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_20_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_20_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_21_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_21_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_21_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_22_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_22_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_22_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_23_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_23_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_23_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_24_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_24_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_24_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_25_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_25_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_25_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_26_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_26_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_26_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_27_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_27_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_27_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_28_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_28_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_28_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_29_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_29_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_29_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_30_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_30_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_30_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_31_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_31_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_31_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_32_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_32_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_32_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_33_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_33_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_33_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_34_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_34_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_34_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_35_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_35_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_35_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_36_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_36_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_36_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_37_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_37_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_37_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_38_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_38_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_38_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_39_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_39_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_39_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_40_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_40_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_40_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_41_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_41_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_41_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_42_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_42_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_42_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_43_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_43_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_43_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_44_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_44_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_44_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_45_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_45_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_45_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_46_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_46_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_46_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_47_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_47_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_47_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_48_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_48_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_48_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_49_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_49_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_49_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_50_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_50_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_50_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_51_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_51_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_51_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_52_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_52_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_52_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_53_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_53_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_53_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_54_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_54_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_54_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_55_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_55_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_55_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_56_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_56_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_56_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_57_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_57_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_57_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_58_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_58_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_58_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_59_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_59_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_59_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_60_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_60_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_60_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_61_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_61_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_61_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_62_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_62_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_62_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_63_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskOut_63_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskOut_63_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_0_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_0_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_0_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_1_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_1_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_1_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_2_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_2_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_2_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_3_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_3_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_3_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_4_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_4_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_4_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_5_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_5_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_5_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_6_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_6_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_6_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_7_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_7_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_7_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_8_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_8_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_8_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_9_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_9_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_9_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_10_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_10_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_10_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_11_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_11_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_11_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_12_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_12_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_12_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_13_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_13_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_13_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_14_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_14_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_14_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_15_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_15_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_15_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_16_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_16_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_16_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_17_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_17_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_17_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_18_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_18_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_18_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_19_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_19_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_19_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_20_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_20_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_20_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_21_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_21_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_21_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_22_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_22_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_22_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_23_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_23_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_23_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_24_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_24_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_24_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_25_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_25_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_25_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_26_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_26_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_26_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_27_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_27_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_27_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_28_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_28_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_28_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_29_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_29_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_29_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_30_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_30_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_30_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_31_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_31_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_31_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_32_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_32_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_32_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_33_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_33_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_33_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_34_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_34_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_34_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_35_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_35_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_35_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_36_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_36_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_36_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_37_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_37_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_37_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_38_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_38_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_38_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_39_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_39_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_39_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_40_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_40_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_40_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_41_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_41_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_41_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_42_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_42_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_42_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_43_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_43_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_43_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_44_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_44_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_44_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_45_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_45_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_45_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_46_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_46_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_46_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_47_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_47_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_47_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_48_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_48_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_48_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_49_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_49_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_49_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_50_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_50_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_50_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_51_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_51_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_51_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_52_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_52_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_52_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_53_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_53_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_53_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_54_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_54_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_54_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_55_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_55_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_55_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_56_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_56_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_56_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_57_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_57_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_57_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_58_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_58_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_58_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_59_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_59_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_59_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_60_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_60_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_60_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_61_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_61_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_61_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_62_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_62_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_62_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_63_TREADY; // @[fullSysGen.scala 228:29]
  wire  stealSide_io_taskIn_63_TVALID; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_io_taskIn_63_TDATA; // @[fullSysGen.scala 228:29]
  wire  stealSide_connSyncSide_0_ctrl_serveStealReq_ready; // @[fullSysGen.scala 228:29]
  wire  stealSide_connSyncSide_0_ctrl_serveStealReq_valid; // @[fullSysGen.scala 228:29]
  wire  stealSide_connSyncSide_0_data_qOutTask_ready; // @[fullSysGen.scala 228:29]
  wire  stealSide_connSyncSide_0_data_qOutTask_valid; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_connSyncSide_0_data_qOutTask_bits; // @[fullSysGen.scala 228:29]
  wire  stealSide_connSyncSide_1_ctrl_serveStealReq_ready; // @[fullSysGen.scala 228:29]
  wire  stealSide_connSyncSide_1_ctrl_serveStealReq_valid; // @[fullSysGen.scala 228:29]
  wire  stealSide_connSyncSide_1_data_qOutTask_ready; // @[fullSysGen.scala 228:29]
  wire  stealSide_connSyncSide_1_data_qOutTask_valid; // @[fullSysGen.scala 228:29]
  wire [255:0] stealSide_connSyncSide_1_data_qOutTask_bits; // @[fullSysGen.scala 228:29]
  wire  continuationAllocationSide_clock; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_reset; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_0_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_0_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_0_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_1_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_1_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_1_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_2_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_2_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_2_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_3_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_3_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_3_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_4_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_4_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_4_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_5_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_5_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_5_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_6_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_6_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_6_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_7_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_7_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_7_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_8_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_8_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_8_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_9_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_9_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_9_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_10_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_10_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_10_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_11_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_11_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_11_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_12_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_12_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_12_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_13_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_13_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_13_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_14_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_14_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_14_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_15_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_15_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_15_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_16_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_16_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_16_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_17_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_17_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_17_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_18_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_18_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_18_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_19_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_19_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_19_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_20_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_20_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_20_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_21_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_21_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_21_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_22_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_22_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_22_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_23_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_23_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_23_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_24_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_24_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_24_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_25_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_25_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_25_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_26_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_26_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_26_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_27_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_27_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_27_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_28_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_28_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_28_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_29_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_29_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_29_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_30_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_30_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_30_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_31_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_31_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_31_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_32_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_32_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_32_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_33_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_33_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_33_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_34_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_34_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_34_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_35_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_35_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_35_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_36_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_36_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_36_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_37_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_37_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_37_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_38_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_38_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_38_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_39_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_39_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_39_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_40_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_40_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_40_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_41_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_41_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_41_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_42_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_42_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_42_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_43_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_43_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_43_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_44_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_44_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_44_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_45_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_45_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_45_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_46_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_46_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_46_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_47_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_47_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_47_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_48_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_48_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_48_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_49_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_49_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_49_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_50_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_50_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_50_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_51_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_51_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_51_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_52_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_52_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_52_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_53_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_53_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_53_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_54_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_54_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_54_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_55_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_55_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_55_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_56_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_56_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_56_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_57_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_57_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_57_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_58_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_58_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_58_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_59_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_59_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_59_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_60_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_60_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_60_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_61_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_61_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_61_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_62_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_62_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_62_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_63_TREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_contOut_63_TVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_contOut_63_TDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_axi_mgmt_vcas_0_ARREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_axi_mgmt_vcas_0_ARVALID; // @[fullSysGen.scala 270:48]
  wire [5:0] continuationAllocationSide_io_axi_mgmt_vcas_0_ARADDR; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_axi_mgmt_vcas_0_RREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_axi_mgmt_vcas_0_RVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_axi_mgmt_vcas_0_RDATA; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_axi_mgmt_vcas_0_AWREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_axi_mgmt_vcas_0_AWVALID; // @[fullSysGen.scala 270:48]
  wire [5:0] continuationAllocationSide_io_axi_mgmt_vcas_0_AWADDR; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_axi_mgmt_vcas_0_WREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_axi_mgmt_vcas_0_WVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_axi_mgmt_vcas_0_WDATA; // @[fullSysGen.scala 270:48]
  wire [7:0] continuationAllocationSide_io_axi_mgmt_vcas_0_WSTRB; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_axi_mgmt_vcas_0_BREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_axi_mgmt_vcas_0_BVALID; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_vcas_axi_full_0_ARREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_vcas_axi_full_0_ARVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_vcas_axi_full_0_ARADDR; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_vcas_axi_full_0_RREADY; // @[fullSysGen.scala 270:48]
  wire  continuationAllocationSide_io_vcas_axi_full_0_RVALID; // @[fullSysGen.scala 270:48]
  wire [63:0] continuationAllocationSide_io_vcas_axi_full_0_RDATA; // @[fullSysGen.scala 270:48]
  wire  syncSide_clock; // @[fullSysGen.scala 284:30]
  wire  syncSide_reset; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_0_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_0_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_0_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_1_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_1_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_1_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_2_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_2_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_2_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_3_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_3_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_3_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_4_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_4_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_4_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_5_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_5_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_5_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_6_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_6_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_6_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_7_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_7_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_7_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_8_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_8_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_8_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_9_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_9_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_9_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_10_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_10_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_10_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_11_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_11_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_11_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_12_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_12_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_12_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_13_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_13_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_13_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_14_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_14_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_14_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_15_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_15_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_15_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_16_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_16_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_16_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_17_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_17_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_17_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_18_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_18_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_18_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_19_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_19_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_19_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_20_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_20_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_20_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_21_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_21_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_21_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_22_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_22_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_22_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_23_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_23_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_23_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_24_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_24_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_24_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_25_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_25_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_25_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_26_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_26_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_26_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_27_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_27_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_27_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_28_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_28_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_28_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_29_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_29_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_29_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_30_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_30_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_30_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_31_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_31_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_31_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_32_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_32_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_32_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_33_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_33_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_33_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_34_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_34_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_34_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_35_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_35_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_35_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_36_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_36_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_36_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_37_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_37_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_37_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_38_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_38_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_38_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_39_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_39_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_39_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_40_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_40_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_40_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_41_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_41_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_41_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_42_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_42_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_42_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_43_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_43_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_43_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_44_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_44_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_44_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_45_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_45_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_45_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_46_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_46_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_46_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_47_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_47_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_47_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_48_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_48_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_48_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_49_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_49_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_49_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_50_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_50_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_50_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_51_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_51_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_51_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_52_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_52_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_52_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_53_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_53_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_53_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_54_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_54_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_54_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_55_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_55_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_55_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_56_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_56_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_56_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_57_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_57_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_57_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_58_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_58_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_58_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_59_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_59_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_59_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_60_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_60_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_60_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_61_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_61_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_61_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_62_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_62_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_62_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_63_TREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_addrIn_63_TVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_addrIn_63_TDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_0_ARREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_0_ARVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_axi_full_argRoute_0_ARADDR; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_0_RREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_0_RVALID; // @[fullSysGen.scala 284:30]
  wire [31:0] syncSide_io_axi_full_argRoute_0_RDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_0_AWREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_0_AWVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_axi_full_argRoute_0_AWADDR; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_0_WREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_0_WVALID; // @[fullSysGen.scala 284:30]
  wire [31:0] syncSide_io_axi_full_argRoute_0_WDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_0_BVALID; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_1_ARREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_1_ARVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_axi_full_argRoute_1_ARADDR; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_1_RREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_1_RVALID; // @[fullSysGen.scala 284:30]
  wire [31:0] syncSide_io_axi_full_argRoute_1_RDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_1_AWREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_1_AWVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_axi_full_argRoute_1_AWADDR; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_1_WREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_1_WVALID; // @[fullSysGen.scala 284:30]
  wire [31:0] syncSide_io_axi_full_argRoute_1_WDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_1_BVALID; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_2_ARREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_2_ARVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_axi_full_argRoute_2_ARADDR; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_2_RREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_2_RVALID; // @[fullSysGen.scala 284:30]
  wire [31:0] syncSide_io_axi_full_argRoute_2_RDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_3_ARREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_3_ARVALID; // @[fullSysGen.scala 284:30]
  wire [63:0] syncSide_io_axi_full_argRoute_3_ARADDR; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_3_RREADY; // @[fullSysGen.scala 284:30]
  wire  syncSide_io_axi_full_argRoute_3_RVALID; // @[fullSysGen.scala 284:30]
  wire [31:0] syncSide_io_axi_full_argRoute_3_RDATA; // @[fullSysGen.scala 284:30]
  wire  syncSide_connStealNtw_0_ctrl_serveStealReq_ready; // @[fullSysGen.scala 284:30]
  wire  syncSide_connStealNtw_0_ctrl_serveStealReq_valid; // @[fullSysGen.scala 284:30]
  wire  syncSide_connStealNtw_0_data_qOutTask_ready; // @[fullSysGen.scala 284:30]
  wire  syncSide_connStealNtw_0_data_qOutTask_valid; // @[fullSysGen.scala 284:30]
  wire [255:0] syncSide_connStealNtw_0_data_qOutTask_bits; // @[fullSysGen.scala 284:30]
  wire  syncSide_connStealNtw_1_ctrl_serveStealReq_ready; // @[fullSysGen.scala 284:30]
  wire  syncSide_connStealNtw_1_ctrl_serveStealReq_valid; // @[fullSysGen.scala 284:30]
  wire  syncSide_connStealNtw_1_data_qOutTask_ready; // @[fullSysGen.scala 284:30]
  wire  syncSide_connStealNtw_1_data_qOutTask_valid; // @[fullSysGen.scala 284:30]
  wire [255:0] syncSide_connStealNtw_1_data_qOutTask_bits; // @[fullSysGen.scala 284:30]
  stealSide stealSide ( // @[fullSysGen.scala 228:29]
    .clock(stealSide_clock),
    .reset(stealSide_reset),
    .io_axi_mgmt_vss_0_ARREADY(stealSide_io_axi_mgmt_vss_0_ARREADY),
    .io_axi_mgmt_vss_0_ARVALID(stealSide_io_axi_mgmt_vss_0_ARVALID),
    .io_axi_mgmt_vss_0_ARADDR(stealSide_io_axi_mgmt_vss_0_ARADDR),
    .io_axi_mgmt_vss_0_RREADY(stealSide_io_axi_mgmt_vss_0_RREADY),
    .io_axi_mgmt_vss_0_RVALID(stealSide_io_axi_mgmt_vss_0_RVALID),
    .io_axi_mgmt_vss_0_RDATA(stealSide_io_axi_mgmt_vss_0_RDATA),
    .io_axi_mgmt_vss_0_AWREADY(stealSide_io_axi_mgmt_vss_0_AWREADY),
    .io_axi_mgmt_vss_0_AWVALID(stealSide_io_axi_mgmt_vss_0_AWVALID),
    .io_axi_mgmt_vss_0_AWADDR(stealSide_io_axi_mgmt_vss_0_AWADDR),
    .io_axi_mgmt_vss_0_WREADY(stealSide_io_axi_mgmt_vss_0_WREADY),
    .io_axi_mgmt_vss_0_WVALID(stealSide_io_axi_mgmt_vss_0_WVALID),
    .io_axi_mgmt_vss_0_WDATA(stealSide_io_axi_mgmt_vss_0_WDATA),
    .io_axi_mgmt_vss_0_WSTRB(stealSide_io_axi_mgmt_vss_0_WSTRB),
    .io_axi_mgmt_vss_0_BREADY(stealSide_io_axi_mgmt_vss_0_BREADY),
    .io_axi_mgmt_vss_0_BVALID(stealSide_io_axi_mgmt_vss_0_BVALID),
    .io_vss_axi_full_0_ARREADY(stealSide_io_vss_axi_full_0_ARREADY),
    .io_vss_axi_full_0_ARVALID(stealSide_io_vss_axi_full_0_ARVALID),
    .io_vss_axi_full_0_ARADDR(stealSide_io_vss_axi_full_0_ARADDR),
    .io_vss_axi_full_0_ARLEN(stealSide_io_vss_axi_full_0_ARLEN),
    .io_vss_axi_full_0_RREADY(stealSide_io_vss_axi_full_0_RREADY),
    .io_vss_axi_full_0_RVALID(stealSide_io_vss_axi_full_0_RVALID),
    .io_vss_axi_full_0_RDATA(stealSide_io_vss_axi_full_0_RDATA),
    .io_vss_axi_full_0_AWREADY(stealSide_io_vss_axi_full_0_AWREADY),
    .io_vss_axi_full_0_AWVALID(stealSide_io_vss_axi_full_0_AWVALID),
    .io_vss_axi_full_0_AWADDR(stealSide_io_vss_axi_full_0_AWADDR),
    .io_vss_axi_full_0_AWLEN(stealSide_io_vss_axi_full_0_AWLEN),
    .io_vss_axi_full_0_WREADY(stealSide_io_vss_axi_full_0_WREADY),
    .io_vss_axi_full_0_WVALID(stealSide_io_vss_axi_full_0_WVALID),
    .io_vss_axi_full_0_WDATA(stealSide_io_vss_axi_full_0_WDATA),
    .io_vss_axi_full_0_WLAST(stealSide_io_vss_axi_full_0_WLAST),
    .io_vss_axi_full_0_BVALID(stealSide_io_vss_axi_full_0_BVALID),
    .io_taskOut_0_TREADY(stealSide_io_taskOut_0_TREADY),
    .io_taskOut_0_TVALID(stealSide_io_taskOut_0_TVALID),
    .io_taskOut_0_TDATA(stealSide_io_taskOut_0_TDATA),
    .io_taskOut_1_TREADY(stealSide_io_taskOut_1_TREADY),
    .io_taskOut_1_TVALID(stealSide_io_taskOut_1_TVALID),
    .io_taskOut_1_TDATA(stealSide_io_taskOut_1_TDATA),
    .io_taskOut_2_TREADY(stealSide_io_taskOut_2_TREADY),
    .io_taskOut_2_TVALID(stealSide_io_taskOut_2_TVALID),
    .io_taskOut_2_TDATA(stealSide_io_taskOut_2_TDATA),
    .io_taskOut_3_TREADY(stealSide_io_taskOut_3_TREADY),
    .io_taskOut_3_TVALID(stealSide_io_taskOut_3_TVALID),
    .io_taskOut_3_TDATA(stealSide_io_taskOut_3_TDATA),
    .io_taskOut_4_TREADY(stealSide_io_taskOut_4_TREADY),
    .io_taskOut_4_TVALID(stealSide_io_taskOut_4_TVALID),
    .io_taskOut_4_TDATA(stealSide_io_taskOut_4_TDATA),
    .io_taskOut_5_TREADY(stealSide_io_taskOut_5_TREADY),
    .io_taskOut_5_TVALID(stealSide_io_taskOut_5_TVALID),
    .io_taskOut_5_TDATA(stealSide_io_taskOut_5_TDATA),
    .io_taskOut_6_TREADY(stealSide_io_taskOut_6_TREADY),
    .io_taskOut_6_TVALID(stealSide_io_taskOut_6_TVALID),
    .io_taskOut_6_TDATA(stealSide_io_taskOut_6_TDATA),
    .io_taskOut_7_TREADY(stealSide_io_taskOut_7_TREADY),
    .io_taskOut_7_TVALID(stealSide_io_taskOut_7_TVALID),
    .io_taskOut_7_TDATA(stealSide_io_taskOut_7_TDATA),
    .io_taskOut_8_TREADY(stealSide_io_taskOut_8_TREADY),
    .io_taskOut_8_TVALID(stealSide_io_taskOut_8_TVALID),
    .io_taskOut_8_TDATA(stealSide_io_taskOut_8_TDATA),
    .io_taskOut_9_TREADY(stealSide_io_taskOut_9_TREADY),
    .io_taskOut_9_TVALID(stealSide_io_taskOut_9_TVALID),
    .io_taskOut_9_TDATA(stealSide_io_taskOut_9_TDATA),
    .io_taskOut_10_TREADY(stealSide_io_taskOut_10_TREADY),
    .io_taskOut_10_TVALID(stealSide_io_taskOut_10_TVALID),
    .io_taskOut_10_TDATA(stealSide_io_taskOut_10_TDATA),
    .io_taskOut_11_TREADY(stealSide_io_taskOut_11_TREADY),
    .io_taskOut_11_TVALID(stealSide_io_taskOut_11_TVALID),
    .io_taskOut_11_TDATA(stealSide_io_taskOut_11_TDATA),
    .io_taskOut_12_TREADY(stealSide_io_taskOut_12_TREADY),
    .io_taskOut_12_TVALID(stealSide_io_taskOut_12_TVALID),
    .io_taskOut_12_TDATA(stealSide_io_taskOut_12_TDATA),
    .io_taskOut_13_TREADY(stealSide_io_taskOut_13_TREADY),
    .io_taskOut_13_TVALID(stealSide_io_taskOut_13_TVALID),
    .io_taskOut_13_TDATA(stealSide_io_taskOut_13_TDATA),
    .io_taskOut_14_TREADY(stealSide_io_taskOut_14_TREADY),
    .io_taskOut_14_TVALID(stealSide_io_taskOut_14_TVALID),
    .io_taskOut_14_TDATA(stealSide_io_taskOut_14_TDATA),
    .io_taskOut_15_TREADY(stealSide_io_taskOut_15_TREADY),
    .io_taskOut_15_TVALID(stealSide_io_taskOut_15_TVALID),
    .io_taskOut_15_TDATA(stealSide_io_taskOut_15_TDATA),
    .io_taskOut_16_TREADY(stealSide_io_taskOut_16_TREADY),
    .io_taskOut_16_TVALID(stealSide_io_taskOut_16_TVALID),
    .io_taskOut_16_TDATA(stealSide_io_taskOut_16_TDATA),
    .io_taskOut_17_TREADY(stealSide_io_taskOut_17_TREADY),
    .io_taskOut_17_TVALID(stealSide_io_taskOut_17_TVALID),
    .io_taskOut_17_TDATA(stealSide_io_taskOut_17_TDATA),
    .io_taskOut_18_TREADY(stealSide_io_taskOut_18_TREADY),
    .io_taskOut_18_TVALID(stealSide_io_taskOut_18_TVALID),
    .io_taskOut_18_TDATA(stealSide_io_taskOut_18_TDATA),
    .io_taskOut_19_TREADY(stealSide_io_taskOut_19_TREADY),
    .io_taskOut_19_TVALID(stealSide_io_taskOut_19_TVALID),
    .io_taskOut_19_TDATA(stealSide_io_taskOut_19_TDATA),
    .io_taskOut_20_TREADY(stealSide_io_taskOut_20_TREADY),
    .io_taskOut_20_TVALID(stealSide_io_taskOut_20_TVALID),
    .io_taskOut_20_TDATA(stealSide_io_taskOut_20_TDATA),
    .io_taskOut_21_TREADY(stealSide_io_taskOut_21_TREADY),
    .io_taskOut_21_TVALID(stealSide_io_taskOut_21_TVALID),
    .io_taskOut_21_TDATA(stealSide_io_taskOut_21_TDATA),
    .io_taskOut_22_TREADY(stealSide_io_taskOut_22_TREADY),
    .io_taskOut_22_TVALID(stealSide_io_taskOut_22_TVALID),
    .io_taskOut_22_TDATA(stealSide_io_taskOut_22_TDATA),
    .io_taskOut_23_TREADY(stealSide_io_taskOut_23_TREADY),
    .io_taskOut_23_TVALID(stealSide_io_taskOut_23_TVALID),
    .io_taskOut_23_TDATA(stealSide_io_taskOut_23_TDATA),
    .io_taskOut_24_TREADY(stealSide_io_taskOut_24_TREADY),
    .io_taskOut_24_TVALID(stealSide_io_taskOut_24_TVALID),
    .io_taskOut_24_TDATA(stealSide_io_taskOut_24_TDATA),
    .io_taskOut_25_TREADY(stealSide_io_taskOut_25_TREADY),
    .io_taskOut_25_TVALID(stealSide_io_taskOut_25_TVALID),
    .io_taskOut_25_TDATA(stealSide_io_taskOut_25_TDATA),
    .io_taskOut_26_TREADY(stealSide_io_taskOut_26_TREADY),
    .io_taskOut_26_TVALID(stealSide_io_taskOut_26_TVALID),
    .io_taskOut_26_TDATA(stealSide_io_taskOut_26_TDATA),
    .io_taskOut_27_TREADY(stealSide_io_taskOut_27_TREADY),
    .io_taskOut_27_TVALID(stealSide_io_taskOut_27_TVALID),
    .io_taskOut_27_TDATA(stealSide_io_taskOut_27_TDATA),
    .io_taskOut_28_TREADY(stealSide_io_taskOut_28_TREADY),
    .io_taskOut_28_TVALID(stealSide_io_taskOut_28_TVALID),
    .io_taskOut_28_TDATA(stealSide_io_taskOut_28_TDATA),
    .io_taskOut_29_TREADY(stealSide_io_taskOut_29_TREADY),
    .io_taskOut_29_TVALID(stealSide_io_taskOut_29_TVALID),
    .io_taskOut_29_TDATA(stealSide_io_taskOut_29_TDATA),
    .io_taskOut_30_TREADY(stealSide_io_taskOut_30_TREADY),
    .io_taskOut_30_TVALID(stealSide_io_taskOut_30_TVALID),
    .io_taskOut_30_TDATA(stealSide_io_taskOut_30_TDATA),
    .io_taskOut_31_TREADY(stealSide_io_taskOut_31_TREADY),
    .io_taskOut_31_TVALID(stealSide_io_taskOut_31_TVALID),
    .io_taskOut_31_TDATA(stealSide_io_taskOut_31_TDATA),
    .io_taskOut_32_TREADY(stealSide_io_taskOut_32_TREADY),
    .io_taskOut_32_TVALID(stealSide_io_taskOut_32_TVALID),
    .io_taskOut_32_TDATA(stealSide_io_taskOut_32_TDATA),
    .io_taskOut_33_TREADY(stealSide_io_taskOut_33_TREADY),
    .io_taskOut_33_TVALID(stealSide_io_taskOut_33_TVALID),
    .io_taskOut_33_TDATA(stealSide_io_taskOut_33_TDATA),
    .io_taskOut_34_TREADY(stealSide_io_taskOut_34_TREADY),
    .io_taskOut_34_TVALID(stealSide_io_taskOut_34_TVALID),
    .io_taskOut_34_TDATA(stealSide_io_taskOut_34_TDATA),
    .io_taskOut_35_TREADY(stealSide_io_taskOut_35_TREADY),
    .io_taskOut_35_TVALID(stealSide_io_taskOut_35_TVALID),
    .io_taskOut_35_TDATA(stealSide_io_taskOut_35_TDATA),
    .io_taskOut_36_TREADY(stealSide_io_taskOut_36_TREADY),
    .io_taskOut_36_TVALID(stealSide_io_taskOut_36_TVALID),
    .io_taskOut_36_TDATA(stealSide_io_taskOut_36_TDATA),
    .io_taskOut_37_TREADY(stealSide_io_taskOut_37_TREADY),
    .io_taskOut_37_TVALID(stealSide_io_taskOut_37_TVALID),
    .io_taskOut_37_TDATA(stealSide_io_taskOut_37_TDATA),
    .io_taskOut_38_TREADY(stealSide_io_taskOut_38_TREADY),
    .io_taskOut_38_TVALID(stealSide_io_taskOut_38_TVALID),
    .io_taskOut_38_TDATA(stealSide_io_taskOut_38_TDATA),
    .io_taskOut_39_TREADY(stealSide_io_taskOut_39_TREADY),
    .io_taskOut_39_TVALID(stealSide_io_taskOut_39_TVALID),
    .io_taskOut_39_TDATA(stealSide_io_taskOut_39_TDATA),
    .io_taskOut_40_TREADY(stealSide_io_taskOut_40_TREADY),
    .io_taskOut_40_TVALID(stealSide_io_taskOut_40_TVALID),
    .io_taskOut_40_TDATA(stealSide_io_taskOut_40_TDATA),
    .io_taskOut_41_TREADY(stealSide_io_taskOut_41_TREADY),
    .io_taskOut_41_TVALID(stealSide_io_taskOut_41_TVALID),
    .io_taskOut_41_TDATA(stealSide_io_taskOut_41_TDATA),
    .io_taskOut_42_TREADY(stealSide_io_taskOut_42_TREADY),
    .io_taskOut_42_TVALID(stealSide_io_taskOut_42_TVALID),
    .io_taskOut_42_TDATA(stealSide_io_taskOut_42_TDATA),
    .io_taskOut_43_TREADY(stealSide_io_taskOut_43_TREADY),
    .io_taskOut_43_TVALID(stealSide_io_taskOut_43_TVALID),
    .io_taskOut_43_TDATA(stealSide_io_taskOut_43_TDATA),
    .io_taskOut_44_TREADY(stealSide_io_taskOut_44_TREADY),
    .io_taskOut_44_TVALID(stealSide_io_taskOut_44_TVALID),
    .io_taskOut_44_TDATA(stealSide_io_taskOut_44_TDATA),
    .io_taskOut_45_TREADY(stealSide_io_taskOut_45_TREADY),
    .io_taskOut_45_TVALID(stealSide_io_taskOut_45_TVALID),
    .io_taskOut_45_TDATA(stealSide_io_taskOut_45_TDATA),
    .io_taskOut_46_TREADY(stealSide_io_taskOut_46_TREADY),
    .io_taskOut_46_TVALID(stealSide_io_taskOut_46_TVALID),
    .io_taskOut_46_TDATA(stealSide_io_taskOut_46_TDATA),
    .io_taskOut_47_TREADY(stealSide_io_taskOut_47_TREADY),
    .io_taskOut_47_TVALID(stealSide_io_taskOut_47_TVALID),
    .io_taskOut_47_TDATA(stealSide_io_taskOut_47_TDATA),
    .io_taskOut_48_TREADY(stealSide_io_taskOut_48_TREADY),
    .io_taskOut_48_TVALID(stealSide_io_taskOut_48_TVALID),
    .io_taskOut_48_TDATA(stealSide_io_taskOut_48_TDATA),
    .io_taskOut_49_TREADY(stealSide_io_taskOut_49_TREADY),
    .io_taskOut_49_TVALID(stealSide_io_taskOut_49_TVALID),
    .io_taskOut_49_TDATA(stealSide_io_taskOut_49_TDATA),
    .io_taskOut_50_TREADY(stealSide_io_taskOut_50_TREADY),
    .io_taskOut_50_TVALID(stealSide_io_taskOut_50_TVALID),
    .io_taskOut_50_TDATA(stealSide_io_taskOut_50_TDATA),
    .io_taskOut_51_TREADY(stealSide_io_taskOut_51_TREADY),
    .io_taskOut_51_TVALID(stealSide_io_taskOut_51_TVALID),
    .io_taskOut_51_TDATA(stealSide_io_taskOut_51_TDATA),
    .io_taskOut_52_TREADY(stealSide_io_taskOut_52_TREADY),
    .io_taskOut_52_TVALID(stealSide_io_taskOut_52_TVALID),
    .io_taskOut_52_TDATA(stealSide_io_taskOut_52_TDATA),
    .io_taskOut_53_TREADY(stealSide_io_taskOut_53_TREADY),
    .io_taskOut_53_TVALID(stealSide_io_taskOut_53_TVALID),
    .io_taskOut_53_TDATA(stealSide_io_taskOut_53_TDATA),
    .io_taskOut_54_TREADY(stealSide_io_taskOut_54_TREADY),
    .io_taskOut_54_TVALID(stealSide_io_taskOut_54_TVALID),
    .io_taskOut_54_TDATA(stealSide_io_taskOut_54_TDATA),
    .io_taskOut_55_TREADY(stealSide_io_taskOut_55_TREADY),
    .io_taskOut_55_TVALID(stealSide_io_taskOut_55_TVALID),
    .io_taskOut_55_TDATA(stealSide_io_taskOut_55_TDATA),
    .io_taskOut_56_TREADY(stealSide_io_taskOut_56_TREADY),
    .io_taskOut_56_TVALID(stealSide_io_taskOut_56_TVALID),
    .io_taskOut_56_TDATA(stealSide_io_taskOut_56_TDATA),
    .io_taskOut_57_TREADY(stealSide_io_taskOut_57_TREADY),
    .io_taskOut_57_TVALID(stealSide_io_taskOut_57_TVALID),
    .io_taskOut_57_TDATA(stealSide_io_taskOut_57_TDATA),
    .io_taskOut_58_TREADY(stealSide_io_taskOut_58_TREADY),
    .io_taskOut_58_TVALID(stealSide_io_taskOut_58_TVALID),
    .io_taskOut_58_TDATA(stealSide_io_taskOut_58_TDATA),
    .io_taskOut_59_TREADY(stealSide_io_taskOut_59_TREADY),
    .io_taskOut_59_TVALID(stealSide_io_taskOut_59_TVALID),
    .io_taskOut_59_TDATA(stealSide_io_taskOut_59_TDATA),
    .io_taskOut_60_TREADY(stealSide_io_taskOut_60_TREADY),
    .io_taskOut_60_TVALID(stealSide_io_taskOut_60_TVALID),
    .io_taskOut_60_TDATA(stealSide_io_taskOut_60_TDATA),
    .io_taskOut_61_TREADY(stealSide_io_taskOut_61_TREADY),
    .io_taskOut_61_TVALID(stealSide_io_taskOut_61_TVALID),
    .io_taskOut_61_TDATA(stealSide_io_taskOut_61_TDATA),
    .io_taskOut_62_TREADY(stealSide_io_taskOut_62_TREADY),
    .io_taskOut_62_TVALID(stealSide_io_taskOut_62_TVALID),
    .io_taskOut_62_TDATA(stealSide_io_taskOut_62_TDATA),
    .io_taskOut_63_TREADY(stealSide_io_taskOut_63_TREADY),
    .io_taskOut_63_TVALID(stealSide_io_taskOut_63_TVALID),
    .io_taskOut_63_TDATA(stealSide_io_taskOut_63_TDATA),
    .io_taskIn_0_TREADY(stealSide_io_taskIn_0_TREADY),
    .io_taskIn_0_TVALID(stealSide_io_taskIn_0_TVALID),
    .io_taskIn_0_TDATA(stealSide_io_taskIn_0_TDATA),
    .io_taskIn_1_TREADY(stealSide_io_taskIn_1_TREADY),
    .io_taskIn_1_TVALID(stealSide_io_taskIn_1_TVALID),
    .io_taskIn_1_TDATA(stealSide_io_taskIn_1_TDATA),
    .io_taskIn_2_TREADY(stealSide_io_taskIn_2_TREADY),
    .io_taskIn_2_TVALID(stealSide_io_taskIn_2_TVALID),
    .io_taskIn_2_TDATA(stealSide_io_taskIn_2_TDATA),
    .io_taskIn_3_TREADY(stealSide_io_taskIn_3_TREADY),
    .io_taskIn_3_TVALID(stealSide_io_taskIn_3_TVALID),
    .io_taskIn_3_TDATA(stealSide_io_taskIn_3_TDATA),
    .io_taskIn_4_TREADY(stealSide_io_taskIn_4_TREADY),
    .io_taskIn_4_TVALID(stealSide_io_taskIn_4_TVALID),
    .io_taskIn_4_TDATA(stealSide_io_taskIn_4_TDATA),
    .io_taskIn_5_TREADY(stealSide_io_taskIn_5_TREADY),
    .io_taskIn_5_TVALID(stealSide_io_taskIn_5_TVALID),
    .io_taskIn_5_TDATA(stealSide_io_taskIn_5_TDATA),
    .io_taskIn_6_TREADY(stealSide_io_taskIn_6_TREADY),
    .io_taskIn_6_TVALID(stealSide_io_taskIn_6_TVALID),
    .io_taskIn_6_TDATA(stealSide_io_taskIn_6_TDATA),
    .io_taskIn_7_TREADY(stealSide_io_taskIn_7_TREADY),
    .io_taskIn_7_TVALID(stealSide_io_taskIn_7_TVALID),
    .io_taskIn_7_TDATA(stealSide_io_taskIn_7_TDATA),
    .io_taskIn_8_TREADY(stealSide_io_taskIn_8_TREADY),
    .io_taskIn_8_TVALID(stealSide_io_taskIn_8_TVALID),
    .io_taskIn_8_TDATA(stealSide_io_taskIn_8_TDATA),
    .io_taskIn_9_TREADY(stealSide_io_taskIn_9_TREADY),
    .io_taskIn_9_TVALID(stealSide_io_taskIn_9_TVALID),
    .io_taskIn_9_TDATA(stealSide_io_taskIn_9_TDATA),
    .io_taskIn_10_TREADY(stealSide_io_taskIn_10_TREADY),
    .io_taskIn_10_TVALID(stealSide_io_taskIn_10_TVALID),
    .io_taskIn_10_TDATA(stealSide_io_taskIn_10_TDATA),
    .io_taskIn_11_TREADY(stealSide_io_taskIn_11_TREADY),
    .io_taskIn_11_TVALID(stealSide_io_taskIn_11_TVALID),
    .io_taskIn_11_TDATA(stealSide_io_taskIn_11_TDATA),
    .io_taskIn_12_TREADY(stealSide_io_taskIn_12_TREADY),
    .io_taskIn_12_TVALID(stealSide_io_taskIn_12_TVALID),
    .io_taskIn_12_TDATA(stealSide_io_taskIn_12_TDATA),
    .io_taskIn_13_TREADY(stealSide_io_taskIn_13_TREADY),
    .io_taskIn_13_TVALID(stealSide_io_taskIn_13_TVALID),
    .io_taskIn_13_TDATA(stealSide_io_taskIn_13_TDATA),
    .io_taskIn_14_TREADY(stealSide_io_taskIn_14_TREADY),
    .io_taskIn_14_TVALID(stealSide_io_taskIn_14_TVALID),
    .io_taskIn_14_TDATA(stealSide_io_taskIn_14_TDATA),
    .io_taskIn_15_TREADY(stealSide_io_taskIn_15_TREADY),
    .io_taskIn_15_TVALID(stealSide_io_taskIn_15_TVALID),
    .io_taskIn_15_TDATA(stealSide_io_taskIn_15_TDATA),
    .io_taskIn_16_TREADY(stealSide_io_taskIn_16_TREADY),
    .io_taskIn_16_TVALID(stealSide_io_taskIn_16_TVALID),
    .io_taskIn_16_TDATA(stealSide_io_taskIn_16_TDATA),
    .io_taskIn_17_TREADY(stealSide_io_taskIn_17_TREADY),
    .io_taskIn_17_TVALID(stealSide_io_taskIn_17_TVALID),
    .io_taskIn_17_TDATA(stealSide_io_taskIn_17_TDATA),
    .io_taskIn_18_TREADY(stealSide_io_taskIn_18_TREADY),
    .io_taskIn_18_TVALID(stealSide_io_taskIn_18_TVALID),
    .io_taskIn_18_TDATA(stealSide_io_taskIn_18_TDATA),
    .io_taskIn_19_TREADY(stealSide_io_taskIn_19_TREADY),
    .io_taskIn_19_TVALID(stealSide_io_taskIn_19_TVALID),
    .io_taskIn_19_TDATA(stealSide_io_taskIn_19_TDATA),
    .io_taskIn_20_TREADY(stealSide_io_taskIn_20_TREADY),
    .io_taskIn_20_TVALID(stealSide_io_taskIn_20_TVALID),
    .io_taskIn_20_TDATA(stealSide_io_taskIn_20_TDATA),
    .io_taskIn_21_TREADY(stealSide_io_taskIn_21_TREADY),
    .io_taskIn_21_TVALID(stealSide_io_taskIn_21_TVALID),
    .io_taskIn_21_TDATA(stealSide_io_taskIn_21_TDATA),
    .io_taskIn_22_TREADY(stealSide_io_taskIn_22_TREADY),
    .io_taskIn_22_TVALID(stealSide_io_taskIn_22_TVALID),
    .io_taskIn_22_TDATA(stealSide_io_taskIn_22_TDATA),
    .io_taskIn_23_TREADY(stealSide_io_taskIn_23_TREADY),
    .io_taskIn_23_TVALID(stealSide_io_taskIn_23_TVALID),
    .io_taskIn_23_TDATA(stealSide_io_taskIn_23_TDATA),
    .io_taskIn_24_TREADY(stealSide_io_taskIn_24_TREADY),
    .io_taskIn_24_TVALID(stealSide_io_taskIn_24_TVALID),
    .io_taskIn_24_TDATA(stealSide_io_taskIn_24_TDATA),
    .io_taskIn_25_TREADY(stealSide_io_taskIn_25_TREADY),
    .io_taskIn_25_TVALID(stealSide_io_taskIn_25_TVALID),
    .io_taskIn_25_TDATA(stealSide_io_taskIn_25_TDATA),
    .io_taskIn_26_TREADY(stealSide_io_taskIn_26_TREADY),
    .io_taskIn_26_TVALID(stealSide_io_taskIn_26_TVALID),
    .io_taskIn_26_TDATA(stealSide_io_taskIn_26_TDATA),
    .io_taskIn_27_TREADY(stealSide_io_taskIn_27_TREADY),
    .io_taskIn_27_TVALID(stealSide_io_taskIn_27_TVALID),
    .io_taskIn_27_TDATA(stealSide_io_taskIn_27_TDATA),
    .io_taskIn_28_TREADY(stealSide_io_taskIn_28_TREADY),
    .io_taskIn_28_TVALID(stealSide_io_taskIn_28_TVALID),
    .io_taskIn_28_TDATA(stealSide_io_taskIn_28_TDATA),
    .io_taskIn_29_TREADY(stealSide_io_taskIn_29_TREADY),
    .io_taskIn_29_TVALID(stealSide_io_taskIn_29_TVALID),
    .io_taskIn_29_TDATA(stealSide_io_taskIn_29_TDATA),
    .io_taskIn_30_TREADY(stealSide_io_taskIn_30_TREADY),
    .io_taskIn_30_TVALID(stealSide_io_taskIn_30_TVALID),
    .io_taskIn_30_TDATA(stealSide_io_taskIn_30_TDATA),
    .io_taskIn_31_TREADY(stealSide_io_taskIn_31_TREADY),
    .io_taskIn_31_TVALID(stealSide_io_taskIn_31_TVALID),
    .io_taskIn_31_TDATA(stealSide_io_taskIn_31_TDATA),
    .io_taskIn_32_TREADY(stealSide_io_taskIn_32_TREADY),
    .io_taskIn_32_TVALID(stealSide_io_taskIn_32_TVALID),
    .io_taskIn_32_TDATA(stealSide_io_taskIn_32_TDATA),
    .io_taskIn_33_TREADY(stealSide_io_taskIn_33_TREADY),
    .io_taskIn_33_TVALID(stealSide_io_taskIn_33_TVALID),
    .io_taskIn_33_TDATA(stealSide_io_taskIn_33_TDATA),
    .io_taskIn_34_TREADY(stealSide_io_taskIn_34_TREADY),
    .io_taskIn_34_TVALID(stealSide_io_taskIn_34_TVALID),
    .io_taskIn_34_TDATA(stealSide_io_taskIn_34_TDATA),
    .io_taskIn_35_TREADY(stealSide_io_taskIn_35_TREADY),
    .io_taskIn_35_TVALID(stealSide_io_taskIn_35_TVALID),
    .io_taskIn_35_TDATA(stealSide_io_taskIn_35_TDATA),
    .io_taskIn_36_TREADY(stealSide_io_taskIn_36_TREADY),
    .io_taskIn_36_TVALID(stealSide_io_taskIn_36_TVALID),
    .io_taskIn_36_TDATA(stealSide_io_taskIn_36_TDATA),
    .io_taskIn_37_TREADY(stealSide_io_taskIn_37_TREADY),
    .io_taskIn_37_TVALID(stealSide_io_taskIn_37_TVALID),
    .io_taskIn_37_TDATA(stealSide_io_taskIn_37_TDATA),
    .io_taskIn_38_TREADY(stealSide_io_taskIn_38_TREADY),
    .io_taskIn_38_TVALID(stealSide_io_taskIn_38_TVALID),
    .io_taskIn_38_TDATA(stealSide_io_taskIn_38_TDATA),
    .io_taskIn_39_TREADY(stealSide_io_taskIn_39_TREADY),
    .io_taskIn_39_TVALID(stealSide_io_taskIn_39_TVALID),
    .io_taskIn_39_TDATA(stealSide_io_taskIn_39_TDATA),
    .io_taskIn_40_TREADY(stealSide_io_taskIn_40_TREADY),
    .io_taskIn_40_TVALID(stealSide_io_taskIn_40_TVALID),
    .io_taskIn_40_TDATA(stealSide_io_taskIn_40_TDATA),
    .io_taskIn_41_TREADY(stealSide_io_taskIn_41_TREADY),
    .io_taskIn_41_TVALID(stealSide_io_taskIn_41_TVALID),
    .io_taskIn_41_TDATA(stealSide_io_taskIn_41_TDATA),
    .io_taskIn_42_TREADY(stealSide_io_taskIn_42_TREADY),
    .io_taskIn_42_TVALID(stealSide_io_taskIn_42_TVALID),
    .io_taskIn_42_TDATA(stealSide_io_taskIn_42_TDATA),
    .io_taskIn_43_TREADY(stealSide_io_taskIn_43_TREADY),
    .io_taskIn_43_TVALID(stealSide_io_taskIn_43_TVALID),
    .io_taskIn_43_TDATA(stealSide_io_taskIn_43_TDATA),
    .io_taskIn_44_TREADY(stealSide_io_taskIn_44_TREADY),
    .io_taskIn_44_TVALID(stealSide_io_taskIn_44_TVALID),
    .io_taskIn_44_TDATA(stealSide_io_taskIn_44_TDATA),
    .io_taskIn_45_TREADY(stealSide_io_taskIn_45_TREADY),
    .io_taskIn_45_TVALID(stealSide_io_taskIn_45_TVALID),
    .io_taskIn_45_TDATA(stealSide_io_taskIn_45_TDATA),
    .io_taskIn_46_TREADY(stealSide_io_taskIn_46_TREADY),
    .io_taskIn_46_TVALID(stealSide_io_taskIn_46_TVALID),
    .io_taskIn_46_TDATA(stealSide_io_taskIn_46_TDATA),
    .io_taskIn_47_TREADY(stealSide_io_taskIn_47_TREADY),
    .io_taskIn_47_TVALID(stealSide_io_taskIn_47_TVALID),
    .io_taskIn_47_TDATA(stealSide_io_taskIn_47_TDATA),
    .io_taskIn_48_TREADY(stealSide_io_taskIn_48_TREADY),
    .io_taskIn_48_TVALID(stealSide_io_taskIn_48_TVALID),
    .io_taskIn_48_TDATA(stealSide_io_taskIn_48_TDATA),
    .io_taskIn_49_TREADY(stealSide_io_taskIn_49_TREADY),
    .io_taskIn_49_TVALID(stealSide_io_taskIn_49_TVALID),
    .io_taskIn_49_TDATA(stealSide_io_taskIn_49_TDATA),
    .io_taskIn_50_TREADY(stealSide_io_taskIn_50_TREADY),
    .io_taskIn_50_TVALID(stealSide_io_taskIn_50_TVALID),
    .io_taskIn_50_TDATA(stealSide_io_taskIn_50_TDATA),
    .io_taskIn_51_TREADY(stealSide_io_taskIn_51_TREADY),
    .io_taskIn_51_TVALID(stealSide_io_taskIn_51_TVALID),
    .io_taskIn_51_TDATA(stealSide_io_taskIn_51_TDATA),
    .io_taskIn_52_TREADY(stealSide_io_taskIn_52_TREADY),
    .io_taskIn_52_TVALID(stealSide_io_taskIn_52_TVALID),
    .io_taskIn_52_TDATA(stealSide_io_taskIn_52_TDATA),
    .io_taskIn_53_TREADY(stealSide_io_taskIn_53_TREADY),
    .io_taskIn_53_TVALID(stealSide_io_taskIn_53_TVALID),
    .io_taskIn_53_TDATA(stealSide_io_taskIn_53_TDATA),
    .io_taskIn_54_TREADY(stealSide_io_taskIn_54_TREADY),
    .io_taskIn_54_TVALID(stealSide_io_taskIn_54_TVALID),
    .io_taskIn_54_TDATA(stealSide_io_taskIn_54_TDATA),
    .io_taskIn_55_TREADY(stealSide_io_taskIn_55_TREADY),
    .io_taskIn_55_TVALID(stealSide_io_taskIn_55_TVALID),
    .io_taskIn_55_TDATA(stealSide_io_taskIn_55_TDATA),
    .io_taskIn_56_TREADY(stealSide_io_taskIn_56_TREADY),
    .io_taskIn_56_TVALID(stealSide_io_taskIn_56_TVALID),
    .io_taskIn_56_TDATA(stealSide_io_taskIn_56_TDATA),
    .io_taskIn_57_TREADY(stealSide_io_taskIn_57_TREADY),
    .io_taskIn_57_TVALID(stealSide_io_taskIn_57_TVALID),
    .io_taskIn_57_TDATA(stealSide_io_taskIn_57_TDATA),
    .io_taskIn_58_TREADY(stealSide_io_taskIn_58_TREADY),
    .io_taskIn_58_TVALID(stealSide_io_taskIn_58_TVALID),
    .io_taskIn_58_TDATA(stealSide_io_taskIn_58_TDATA),
    .io_taskIn_59_TREADY(stealSide_io_taskIn_59_TREADY),
    .io_taskIn_59_TVALID(stealSide_io_taskIn_59_TVALID),
    .io_taskIn_59_TDATA(stealSide_io_taskIn_59_TDATA),
    .io_taskIn_60_TREADY(stealSide_io_taskIn_60_TREADY),
    .io_taskIn_60_TVALID(stealSide_io_taskIn_60_TVALID),
    .io_taskIn_60_TDATA(stealSide_io_taskIn_60_TDATA),
    .io_taskIn_61_TREADY(stealSide_io_taskIn_61_TREADY),
    .io_taskIn_61_TVALID(stealSide_io_taskIn_61_TVALID),
    .io_taskIn_61_TDATA(stealSide_io_taskIn_61_TDATA),
    .io_taskIn_62_TREADY(stealSide_io_taskIn_62_TREADY),
    .io_taskIn_62_TVALID(stealSide_io_taskIn_62_TVALID),
    .io_taskIn_62_TDATA(stealSide_io_taskIn_62_TDATA),
    .io_taskIn_63_TREADY(stealSide_io_taskIn_63_TREADY),
    .io_taskIn_63_TVALID(stealSide_io_taskIn_63_TVALID),
    .io_taskIn_63_TDATA(stealSide_io_taskIn_63_TDATA),
    .connSyncSide_0_ctrl_serveStealReq_ready(stealSide_connSyncSide_0_ctrl_serveStealReq_ready),
    .connSyncSide_0_ctrl_serveStealReq_valid(stealSide_connSyncSide_0_ctrl_serveStealReq_valid),
    .connSyncSide_0_data_qOutTask_ready(stealSide_connSyncSide_0_data_qOutTask_ready),
    .connSyncSide_0_data_qOutTask_valid(stealSide_connSyncSide_0_data_qOutTask_valid),
    .connSyncSide_0_data_qOutTask_bits(stealSide_connSyncSide_0_data_qOutTask_bits),
    .connSyncSide_1_ctrl_serveStealReq_ready(stealSide_connSyncSide_1_ctrl_serveStealReq_ready),
    .connSyncSide_1_ctrl_serveStealReq_valid(stealSide_connSyncSide_1_ctrl_serveStealReq_valid),
    .connSyncSide_1_data_qOutTask_ready(stealSide_connSyncSide_1_data_qOutTask_ready),
    .connSyncSide_1_data_qOutTask_valid(stealSide_connSyncSide_1_data_qOutTask_valid),
    .connSyncSide_1_data_qOutTask_bits(stealSide_connSyncSide_1_data_qOutTask_bits)
  );
  continuationAllocationSide continuationAllocationSide ( // @[fullSysGen.scala 270:48]
    .clock(continuationAllocationSide_clock),
    .reset(continuationAllocationSide_reset),
    .io_contOut_0_TREADY(continuationAllocationSide_io_contOut_0_TREADY),
    .io_contOut_0_TVALID(continuationAllocationSide_io_contOut_0_TVALID),
    .io_contOut_0_TDATA(continuationAllocationSide_io_contOut_0_TDATA),
    .io_contOut_1_TREADY(continuationAllocationSide_io_contOut_1_TREADY),
    .io_contOut_1_TVALID(continuationAllocationSide_io_contOut_1_TVALID),
    .io_contOut_1_TDATA(continuationAllocationSide_io_contOut_1_TDATA),
    .io_contOut_2_TREADY(continuationAllocationSide_io_contOut_2_TREADY),
    .io_contOut_2_TVALID(continuationAllocationSide_io_contOut_2_TVALID),
    .io_contOut_2_TDATA(continuationAllocationSide_io_contOut_2_TDATA),
    .io_contOut_3_TREADY(continuationAllocationSide_io_contOut_3_TREADY),
    .io_contOut_3_TVALID(continuationAllocationSide_io_contOut_3_TVALID),
    .io_contOut_3_TDATA(continuationAllocationSide_io_contOut_3_TDATA),
    .io_contOut_4_TREADY(continuationAllocationSide_io_contOut_4_TREADY),
    .io_contOut_4_TVALID(continuationAllocationSide_io_contOut_4_TVALID),
    .io_contOut_4_TDATA(continuationAllocationSide_io_contOut_4_TDATA),
    .io_contOut_5_TREADY(continuationAllocationSide_io_contOut_5_TREADY),
    .io_contOut_5_TVALID(continuationAllocationSide_io_contOut_5_TVALID),
    .io_contOut_5_TDATA(continuationAllocationSide_io_contOut_5_TDATA),
    .io_contOut_6_TREADY(continuationAllocationSide_io_contOut_6_TREADY),
    .io_contOut_6_TVALID(continuationAllocationSide_io_contOut_6_TVALID),
    .io_contOut_6_TDATA(continuationAllocationSide_io_contOut_6_TDATA),
    .io_contOut_7_TREADY(continuationAllocationSide_io_contOut_7_TREADY),
    .io_contOut_7_TVALID(continuationAllocationSide_io_contOut_7_TVALID),
    .io_contOut_7_TDATA(continuationAllocationSide_io_contOut_7_TDATA),
    .io_contOut_8_TREADY(continuationAllocationSide_io_contOut_8_TREADY),
    .io_contOut_8_TVALID(continuationAllocationSide_io_contOut_8_TVALID),
    .io_contOut_8_TDATA(continuationAllocationSide_io_contOut_8_TDATA),
    .io_contOut_9_TREADY(continuationAllocationSide_io_contOut_9_TREADY),
    .io_contOut_9_TVALID(continuationAllocationSide_io_contOut_9_TVALID),
    .io_contOut_9_TDATA(continuationAllocationSide_io_contOut_9_TDATA),
    .io_contOut_10_TREADY(continuationAllocationSide_io_contOut_10_TREADY),
    .io_contOut_10_TVALID(continuationAllocationSide_io_contOut_10_TVALID),
    .io_contOut_10_TDATA(continuationAllocationSide_io_contOut_10_TDATA),
    .io_contOut_11_TREADY(continuationAllocationSide_io_contOut_11_TREADY),
    .io_contOut_11_TVALID(continuationAllocationSide_io_contOut_11_TVALID),
    .io_contOut_11_TDATA(continuationAllocationSide_io_contOut_11_TDATA),
    .io_contOut_12_TREADY(continuationAllocationSide_io_contOut_12_TREADY),
    .io_contOut_12_TVALID(continuationAllocationSide_io_contOut_12_TVALID),
    .io_contOut_12_TDATA(continuationAllocationSide_io_contOut_12_TDATA),
    .io_contOut_13_TREADY(continuationAllocationSide_io_contOut_13_TREADY),
    .io_contOut_13_TVALID(continuationAllocationSide_io_contOut_13_TVALID),
    .io_contOut_13_TDATA(continuationAllocationSide_io_contOut_13_TDATA),
    .io_contOut_14_TREADY(continuationAllocationSide_io_contOut_14_TREADY),
    .io_contOut_14_TVALID(continuationAllocationSide_io_contOut_14_TVALID),
    .io_contOut_14_TDATA(continuationAllocationSide_io_contOut_14_TDATA),
    .io_contOut_15_TREADY(continuationAllocationSide_io_contOut_15_TREADY),
    .io_contOut_15_TVALID(continuationAllocationSide_io_contOut_15_TVALID),
    .io_contOut_15_TDATA(continuationAllocationSide_io_contOut_15_TDATA),
    .io_contOut_16_TREADY(continuationAllocationSide_io_contOut_16_TREADY),
    .io_contOut_16_TVALID(continuationAllocationSide_io_contOut_16_TVALID),
    .io_contOut_16_TDATA(continuationAllocationSide_io_contOut_16_TDATA),
    .io_contOut_17_TREADY(continuationAllocationSide_io_contOut_17_TREADY),
    .io_contOut_17_TVALID(continuationAllocationSide_io_contOut_17_TVALID),
    .io_contOut_17_TDATA(continuationAllocationSide_io_contOut_17_TDATA),
    .io_contOut_18_TREADY(continuationAllocationSide_io_contOut_18_TREADY),
    .io_contOut_18_TVALID(continuationAllocationSide_io_contOut_18_TVALID),
    .io_contOut_18_TDATA(continuationAllocationSide_io_contOut_18_TDATA),
    .io_contOut_19_TREADY(continuationAllocationSide_io_contOut_19_TREADY),
    .io_contOut_19_TVALID(continuationAllocationSide_io_contOut_19_TVALID),
    .io_contOut_19_TDATA(continuationAllocationSide_io_contOut_19_TDATA),
    .io_contOut_20_TREADY(continuationAllocationSide_io_contOut_20_TREADY),
    .io_contOut_20_TVALID(continuationAllocationSide_io_contOut_20_TVALID),
    .io_contOut_20_TDATA(continuationAllocationSide_io_contOut_20_TDATA),
    .io_contOut_21_TREADY(continuationAllocationSide_io_contOut_21_TREADY),
    .io_contOut_21_TVALID(continuationAllocationSide_io_contOut_21_TVALID),
    .io_contOut_21_TDATA(continuationAllocationSide_io_contOut_21_TDATA),
    .io_contOut_22_TREADY(continuationAllocationSide_io_contOut_22_TREADY),
    .io_contOut_22_TVALID(continuationAllocationSide_io_contOut_22_TVALID),
    .io_contOut_22_TDATA(continuationAllocationSide_io_contOut_22_TDATA),
    .io_contOut_23_TREADY(continuationAllocationSide_io_contOut_23_TREADY),
    .io_contOut_23_TVALID(continuationAllocationSide_io_contOut_23_TVALID),
    .io_contOut_23_TDATA(continuationAllocationSide_io_contOut_23_TDATA),
    .io_contOut_24_TREADY(continuationAllocationSide_io_contOut_24_TREADY),
    .io_contOut_24_TVALID(continuationAllocationSide_io_contOut_24_TVALID),
    .io_contOut_24_TDATA(continuationAllocationSide_io_contOut_24_TDATA),
    .io_contOut_25_TREADY(continuationAllocationSide_io_contOut_25_TREADY),
    .io_contOut_25_TVALID(continuationAllocationSide_io_contOut_25_TVALID),
    .io_contOut_25_TDATA(continuationAllocationSide_io_contOut_25_TDATA),
    .io_contOut_26_TREADY(continuationAllocationSide_io_contOut_26_TREADY),
    .io_contOut_26_TVALID(continuationAllocationSide_io_contOut_26_TVALID),
    .io_contOut_26_TDATA(continuationAllocationSide_io_contOut_26_TDATA),
    .io_contOut_27_TREADY(continuationAllocationSide_io_contOut_27_TREADY),
    .io_contOut_27_TVALID(continuationAllocationSide_io_contOut_27_TVALID),
    .io_contOut_27_TDATA(continuationAllocationSide_io_contOut_27_TDATA),
    .io_contOut_28_TREADY(continuationAllocationSide_io_contOut_28_TREADY),
    .io_contOut_28_TVALID(continuationAllocationSide_io_contOut_28_TVALID),
    .io_contOut_28_TDATA(continuationAllocationSide_io_contOut_28_TDATA),
    .io_contOut_29_TREADY(continuationAllocationSide_io_contOut_29_TREADY),
    .io_contOut_29_TVALID(continuationAllocationSide_io_contOut_29_TVALID),
    .io_contOut_29_TDATA(continuationAllocationSide_io_contOut_29_TDATA),
    .io_contOut_30_TREADY(continuationAllocationSide_io_contOut_30_TREADY),
    .io_contOut_30_TVALID(continuationAllocationSide_io_contOut_30_TVALID),
    .io_contOut_30_TDATA(continuationAllocationSide_io_contOut_30_TDATA),
    .io_contOut_31_TREADY(continuationAllocationSide_io_contOut_31_TREADY),
    .io_contOut_31_TVALID(continuationAllocationSide_io_contOut_31_TVALID),
    .io_contOut_31_TDATA(continuationAllocationSide_io_contOut_31_TDATA),
    .io_contOut_32_TREADY(continuationAllocationSide_io_contOut_32_TREADY),
    .io_contOut_32_TVALID(continuationAllocationSide_io_contOut_32_TVALID),
    .io_contOut_32_TDATA(continuationAllocationSide_io_contOut_32_TDATA),
    .io_contOut_33_TREADY(continuationAllocationSide_io_contOut_33_TREADY),
    .io_contOut_33_TVALID(continuationAllocationSide_io_contOut_33_TVALID),
    .io_contOut_33_TDATA(continuationAllocationSide_io_contOut_33_TDATA),
    .io_contOut_34_TREADY(continuationAllocationSide_io_contOut_34_TREADY),
    .io_contOut_34_TVALID(continuationAllocationSide_io_contOut_34_TVALID),
    .io_contOut_34_TDATA(continuationAllocationSide_io_contOut_34_TDATA),
    .io_contOut_35_TREADY(continuationAllocationSide_io_contOut_35_TREADY),
    .io_contOut_35_TVALID(continuationAllocationSide_io_contOut_35_TVALID),
    .io_contOut_35_TDATA(continuationAllocationSide_io_contOut_35_TDATA),
    .io_contOut_36_TREADY(continuationAllocationSide_io_contOut_36_TREADY),
    .io_contOut_36_TVALID(continuationAllocationSide_io_contOut_36_TVALID),
    .io_contOut_36_TDATA(continuationAllocationSide_io_contOut_36_TDATA),
    .io_contOut_37_TREADY(continuationAllocationSide_io_contOut_37_TREADY),
    .io_contOut_37_TVALID(continuationAllocationSide_io_contOut_37_TVALID),
    .io_contOut_37_TDATA(continuationAllocationSide_io_contOut_37_TDATA),
    .io_contOut_38_TREADY(continuationAllocationSide_io_contOut_38_TREADY),
    .io_contOut_38_TVALID(continuationAllocationSide_io_contOut_38_TVALID),
    .io_contOut_38_TDATA(continuationAllocationSide_io_contOut_38_TDATA),
    .io_contOut_39_TREADY(continuationAllocationSide_io_contOut_39_TREADY),
    .io_contOut_39_TVALID(continuationAllocationSide_io_contOut_39_TVALID),
    .io_contOut_39_TDATA(continuationAllocationSide_io_contOut_39_TDATA),
    .io_contOut_40_TREADY(continuationAllocationSide_io_contOut_40_TREADY),
    .io_contOut_40_TVALID(continuationAllocationSide_io_contOut_40_TVALID),
    .io_contOut_40_TDATA(continuationAllocationSide_io_contOut_40_TDATA),
    .io_contOut_41_TREADY(continuationAllocationSide_io_contOut_41_TREADY),
    .io_contOut_41_TVALID(continuationAllocationSide_io_contOut_41_TVALID),
    .io_contOut_41_TDATA(continuationAllocationSide_io_contOut_41_TDATA),
    .io_contOut_42_TREADY(continuationAllocationSide_io_contOut_42_TREADY),
    .io_contOut_42_TVALID(continuationAllocationSide_io_contOut_42_TVALID),
    .io_contOut_42_TDATA(continuationAllocationSide_io_contOut_42_TDATA),
    .io_contOut_43_TREADY(continuationAllocationSide_io_contOut_43_TREADY),
    .io_contOut_43_TVALID(continuationAllocationSide_io_contOut_43_TVALID),
    .io_contOut_43_TDATA(continuationAllocationSide_io_contOut_43_TDATA),
    .io_contOut_44_TREADY(continuationAllocationSide_io_contOut_44_TREADY),
    .io_contOut_44_TVALID(continuationAllocationSide_io_contOut_44_TVALID),
    .io_contOut_44_TDATA(continuationAllocationSide_io_contOut_44_TDATA),
    .io_contOut_45_TREADY(continuationAllocationSide_io_contOut_45_TREADY),
    .io_contOut_45_TVALID(continuationAllocationSide_io_contOut_45_TVALID),
    .io_contOut_45_TDATA(continuationAllocationSide_io_contOut_45_TDATA),
    .io_contOut_46_TREADY(continuationAllocationSide_io_contOut_46_TREADY),
    .io_contOut_46_TVALID(continuationAllocationSide_io_contOut_46_TVALID),
    .io_contOut_46_TDATA(continuationAllocationSide_io_contOut_46_TDATA),
    .io_contOut_47_TREADY(continuationAllocationSide_io_contOut_47_TREADY),
    .io_contOut_47_TVALID(continuationAllocationSide_io_contOut_47_TVALID),
    .io_contOut_47_TDATA(continuationAllocationSide_io_contOut_47_TDATA),
    .io_contOut_48_TREADY(continuationAllocationSide_io_contOut_48_TREADY),
    .io_contOut_48_TVALID(continuationAllocationSide_io_contOut_48_TVALID),
    .io_contOut_48_TDATA(continuationAllocationSide_io_contOut_48_TDATA),
    .io_contOut_49_TREADY(continuationAllocationSide_io_contOut_49_TREADY),
    .io_contOut_49_TVALID(continuationAllocationSide_io_contOut_49_TVALID),
    .io_contOut_49_TDATA(continuationAllocationSide_io_contOut_49_TDATA),
    .io_contOut_50_TREADY(continuationAllocationSide_io_contOut_50_TREADY),
    .io_contOut_50_TVALID(continuationAllocationSide_io_contOut_50_TVALID),
    .io_contOut_50_TDATA(continuationAllocationSide_io_contOut_50_TDATA),
    .io_contOut_51_TREADY(continuationAllocationSide_io_contOut_51_TREADY),
    .io_contOut_51_TVALID(continuationAllocationSide_io_contOut_51_TVALID),
    .io_contOut_51_TDATA(continuationAllocationSide_io_contOut_51_TDATA),
    .io_contOut_52_TREADY(continuationAllocationSide_io_contOut_52_TREADY),
    .io_contOut_52_TVALID(continuationAllocationSide_io_contOut_52_TVALID),
    .io_contOut_52_TDATA(continuationAllocationSide_io_contOut_52_TDATA),
    .io_contOut_53_TREADY(continuationAllocationSide_io_contOut_53_TREADY),
    .io_contOut_53_TVALID(continuationAllocationSide_io_contOut_53_TVALID),
    .io_contOut_53_TDATA(continuationAllocationSide_io_contOut_53_TDATA),
    .io_contOut_54_TREADY(continuationAllocationSide_io_contOut_54_TREADY),
    .io_contOut_54_TVALID(continuationAllocationSide_io_contOut_54_TVALID),
    .io_contOut_54_TDATA(continuationAllocationSide_io_contOut_54_TDATA),
    .io_contOut_55_TREADY(continuationAllocationSide_io_contOut_55_TREADY),
    .io_contOut_55_TVALID(continuationAllocationSide_io_contOut_55_TVALID),
    .io_contOut_55_TDATA(continuationAllocationSide_io_contOut_55_TDATA),
    .io_contOut_56_TREADY(continuationAllocationSide_io_contOut_56_TREADY),
    .io_contOut_56_TVALID(continuationAllocationSide_io_contOut_56_TVALID),
    .io_contOut_56_TDATA(continuationAllocationSide_io_contOut_56_TDATA),
    .io_contOut_57_TREADY(continuationAllocationSide_io_contOut_57_TREADY),
    .io_contOut_57_TVALID(continuationAllocationSide_io_contOut_57_TVALID),
    .io_contOut_57_TDATA(continuationAllocationSide_io_contOut_57_TDATA),
    .io_contOut_58_TREADY(continuationAllocationSide_io_contOut_58_TREADY),
    .io_contOut_58_TVALID(continuationAllocationSide_io_contOut_58_TVALID),
    .io_contOut_58_TDATA(continuationAllocationSide_io_contOut_58_TDATA),
    .io_contOut_59_TREADY(continuationAllocationSide_io_contOut_59_TREADY),
    .io_contOut_59_TVALID(continuationAllocationSide_io_contOut_59_TVALID),
    .io_contOut_59_TDATA(continuationAllocationSide_io_contOut_59_TDATA),
    .io_contOut_60_TREADY(continuationAllocationSide_io_contOut_60_TREADY),
    .io_contOut_60_TVALID(continuationAllocationSide_io_contOut_60_TVALID),
    .io_contOut_60_TDATA(continuationAllocationSide_io_contOut_60_TDATA),
    .io_contOut_61_TREADY(continuationAllocationSide_io_contOut_61_TREADY),
    .io_contOut_61_TVALID(continuationAllocationSide_io_contOut_61_TVALID),
    .io_contOut_61_TDATA(continuationAllocationSide_io_contOut_61_TDATA),
    .io_contOut_62_TREADY(continuationAllocationSide_io_contOut_62_TREADY),
    .io_contOut_62_TVALID(continuationAllocationSide_io_contOut_62_TVALID),
    .io_contOut_62_TDATA(continuationAllocationSide_io_contOut_62_TDATA),
    .io_contOut_63_TREADY(continuationAllocationSide_io_contOut_63_TREADY),
    .io_contOut_63_TVALID(continuationAllocationSide_io_contOut_63_TVALID),
    .io_contOut_63_TDATA(continuationAllocationSide_io_contOut_63_TDATA),
    .io_axi_mgmt_vcas_0_ARREADY(continuationAllocationSide_io_axi_mgmt_vcas_0_ARREADY),
    .io_axi_mgmt_vcas_0_ARVALID(continuationAllocationSide_io_axi_mgmt_vcas_0_ARVALID),
    .io_axi_mgmt_vcas_0_ARADDR(continuationAllocationSide_io_axi_mgmt_vcas_0_ARADDR),
    .io_axi_mgmt_vcas_0_RREADY(continuationAllocationSide_io_axi_mgmt_vcas_0_RREADY),
    .io_axi_mgmt_vcas_0_RVALID(continuationAllocationSide_io_axi_mgmt_vcas_0_RVALID),
    .io_axi_mgmt_vcas_0_RDATA(continuationAllocationSide_io_axi_mgmt_vcas_0_RDATA),
    .io_axi_mgmt_vcas_0_AWREADY(continuationAllocationSide_io_axi_mgmt_vcas_0_AWREADY),
    .io_axi_mgmt_vcas_0_AWVALID(continuationAllocationSide_io_axi_mgmt_vcas_0_AWVALID),
    .io_axi_mgmt_vcas_0_AWADDR(continuationAllocationSide_io_axi_mgmt_vcas_0_AWADDR),
    .io_axi_mgmt_vcas_0_WREADY(continuationAllocationSide_io_axi_mgmt_vcas_0_WREADY),
    .io_axi_mgmt_vcas_0_WVALID(continuationAllocationSide_io_axi_mgmt_vcas_0_WVALID),
    .io_axi_mgmt_vcas_0_WDATA(continuationAllocationSide_io_axi_mgmt_vcas_0_WDATA),
    .io_axi_mgmt_vcas_0_WSTRB(continuationAllocationSide_io_axi_mgmt_vcas_0_WSTRB),
    .io_axi_mgmt_vcas_0_BREADY(continuationAllocationSide_io_axi_mgmt_vcas_0_BREADY),
    .io_axi_mgmt_vcas_0_BVALID(continuationAllocationSide_io_axi_mgmt_vcas_0_BVALID),
    .io_vcas_axi_full_0_ARREADY(continuationAllocationSide_io_vcas_axi_full_0_ARREADY),
    .io_vcas_axi_full_0_ARVALID(continuationAllocationSide_io_vcas_axi_full_0_ARVALID),
    .io_vcas_axi_full_0_ARADDR(continuationAllocationSide_io_vcas_axi_full_0_ARADDR),
    .io_vcas_axi_full_0_RREADY(continuationAllocationSide_io_vcas_axi_full_0_RREADY),
    .io_vcas_axi_full_0_RVALID(continuationAllocationSide_io_vcas_axi_full_0_RVALID),
    .io_vcas_axi_full_0_RDATA(continuationAllocationSide_io_vcas_axi_full_0_RDATA)
  );
  syncSide syncSide ( // @[fullSysGen.scala 284:30]
    .clock(syncSide_clock),
    .reset(syncSide_reset),
    .io_addrIn_0_TREADY(syncSide_io_addrIn_0_TREADY),
    .io_addrIn_0_TVALID(syncSide_io_addrIn_0_TVALID),
    .io_addrIn_0_TDATA(syncSide_io_addrIn_0_TDATA),
    .io_addrIn_1_TREADY(syncSide_io_addrIn_1_TREADY),
    .io_addrIn_1_TVALID(syncSide_io_addrIn_1_TVALID),
    .io_addrIn_1_TDATA(syncSide_io_addrIn_1_TDATA),
    .io_addrIn_2_TREADY(syncSide_io_addrIn_2_TREADY),
    .io_addrIn_2_TVALID(syncSide_io_addrIn_2_TVALID),
    .io_addrIn_2_TDATA(syncSide_io_addrIn_2_TDATA),
    .io_addrIn_3_TREADY(syncSide_io_addrIn_3_TREADY),
    .io_addrIn_3_TVALID(syncSide_io_addrIn_3_TVALID),
    .io_addrIn_3_TDATA(syncSide_io_addrIn_3_TDATA),
    .io_addrIn_4_TREADY(syncSide_io_addrIn_4_TREADY),
    .io_addrIn_4_TVALID(syncSide_io_addrIn_4_TVALID),
    .io_addrIn_4_TDATA(syncSide_io_addrIn_4_TDATA),
    .io_addrIn_5_TREADY(syncSide_io_addrIn_5_TREADY),
    .io_addrIn_5_TVALID(syncSide_io_addrIn_5_TVALID),
    .io_addrIn_5_TDATA(syncSide_io_addrIn_5_TDATA),
    .io_addrIn_6_TREADY(syncSide_io_addrIn_6_TREADY),
    .io_addrIn_6_TVALID(syncSide_io_addrIn_6_TVALID),
    .io_addrIn_6_TDATA(syncSide_io_addrIn_6_TDATA),
    .io_addrIn_7_TREADY(syncSide_io_addrIn_7_TREADY),
    .io_addrIn_7_TVALID(syncSide_io_addrIn_7_TVALID),
    .io_addrIn_7_TDATA(syncSide_io_addrIn_7_TDATA),
    .io_addrIn_8_TREADY(syncSide_io_addrIn_8_TREADY),
    .io_addrIn_8_TVALID(syncSide_io_addrIn_8_TVALID),
    .io_addrIn_8_TDATA(syncSide_io_addrIn_8_TDATA),
    .io_addrIn_9_TREADY(syncSide_io_addrIn_9_TREADY),
    .io_addrIn_9_TVALID(syncSide_io_addrIn_9_TVALID),
    .io_addrIn_9_TDATA(syncSide_io_addrIn_9_TDATA),
    .io_addrIn_10_TREADY(syncSide_io_addrIn_10_TREADY),
    .io_addrIn_10_TVALID(syncSide_io_addrIn_10_TVALID),
    .io_addrIn_10_TDATA(syncSide_io_addrIn_10_TDATA),
    .io_addrIn_11_TREADY(syncSide_io_addrIn_11_TREADY),
    .io_addrIn_11_TVALID(syncSide_io_addrIn_11_TVALID),
    .io_addrIn_11_TDATA(syncSide_io_addrIn_11_TDATA),
    .io_addrIn_12_TREADY(syncSide_io_addrIn_12_TREADY),
    .io_addrIn_12_TVALID(syncSide_io_addrIn_12_TVALID),
    .io_addrIn_12_TDATA(syncSide_io_addrIn_12_TDATA),
    .io_addrIn_13_TREADY(syncSide_io_addrIn_13_TREADY),
    .io_addrIn_13_TVALID(syncSide_io_addrIn_13_TVALID),
    .io_addrIn_13_TDATA(syncSide_io_addrIn_13_TDATA),
    .io_addrIn_14_TREADY(syncSide_io_addrIn_14_TREADY),
    .io_addrIn_14_TVALID(syncSide_io_addrIn_14_TVALID),
    .io_addrIn_14_TDATA(syncSide_io_addrIn_14_TDATA),
    .io_addrIn_15_TREADY(syncSide_io_addrIn_15_TREADY),
    .io_addrIn_15_TVALID(syncSide_io_addrIn_15_TVALID),
    .io_addrIn_15_TDATA(syncSide_io_addrIn_15_TDATA),
    .io_addrIn_16_TREADY(syncSide_io_addrIn_16_TREADY),
    .io_addrIn_16_TVALID(syncSide_io_addrIn_16_TVALID),
    .io_addrIn_16_TDATA(syncSide_io_addrIn_16_TDATA),
    .io_addrIn_17_TREADY(syncSide_io_addrIn_17_TREADY),
    .io_addrIn_17_TVALID(syncSide_io_addrIn_17_TVALID),
    .io_addrIn_17_TDATA(syncSide_io_addrIn_17_TDATA),
    .io_addrIn_18_TREADY(syncSide_io_addrIn_18_TREADY),
    .io_addrIn_18_TVALID(syncSide_io_addrIn_18_TVALID),
    .io_addrIn_18_TDATA(syncSide_io_addrIn_18_TDATA),
    .io_addrIn_19_TREADY(syncSide_io_addrIn_19_TREADY),
    .io_addrIn_19_TVALID(syncSide_io_addrIn_19_TVALID),
    .io_addrIn_19_TDATA(syncSide_io_addrIn_19_TDATA),
    .io_addrIn_20_TREADY(syncSide_io_addrIn_20_TREADY),
    .io_addrIn_20_TVALID(syncSide_io_addrIn_20_TVALID),
    .io_addrIn_20_TDATA(syncSide_io_addrIn_20_TDATA),
    .io_addrIn_21_TREADY(syncSide_io_addrIn_21_TREADY),
    .io_addrIn_21_TVALID(syncSide_io_addrIn_21_TVALID),
    .io_addrIn_21_TDATA(syncSide_io_addrIn_21_TDATA),
    .io_addrIn_22_TREADY(syncSide_io_addrIn_22_TREADY),
    .io_addrIn_22_TVALID(syncSide_io_addrIn_22_TVALID),
    .io_addrIn_22_TDATA(syncSide_io_addrIn_22_TDATA),
    .io_addrIn_23_TREADY(syncSide_io_addrIn_23_TREADY),
    .io_addrIn_23_TVALID(syncSide_io_addrIn_23_TVALID),
    .io_addrIn_23_TDATA(syncSide_io_addrIn_23_TDATA),
    .io_addrIn_24_TREADY(syncSide_io_addrIn_24_TREADY),
    .io_addrIn_24_TVALID(syncSide_io_addrIn_24_TVALID),
    .io_addrIn_24_TDATA(syncSide_io_addrIn_24_TDATA),
    .io_addrIn_25_TREADY(syncSide_io_addrIn_25_TREADY),
    .io_addrIn_25_TVALID(syncSide_io_addrIn_25_TVALID),
    .io_addrIn_25_TDATA(syncSide_io_addrIn_25_TDATA),
    .io_addrIn_26_TREADY(syncSide_io_addrIn_26_TREADY),
    .io_addrIn_26_TVALID(syncSide_io_addrIn_26_TVALID),
    .io_addrIn_26_TDATA(syncSide_io_addrIn_26_TDATA),
    .io_addrIn_27_TREADY(syncSide_io_addrIn_27_TREADY),
    .io_addrIn_27_TVALID(syncSide_io_addrIn_27_TVALID),
    .io_addrIn_27_TDATA(syncSide_io_addrIn_27_TDATA),
    .io_addrIn_28_TREADY(syncSide_io_addrIn_28_TREADY),
    .io_addrIn_28_TVALID(syncSide_io_addrIn_28_TVALID),
    .io_addrIn_28_TDATA(syncSide_io_addrIn_28_TDATA),
    .io_addrIn_29_TREADY(syncSide_io_addrIn_29_TREADY),
    .io_addrIn_29_TVALID(syncSide_io_addrIn_29_TVALID),
    .io_addrIn_29_TDATA(syncSide_io_addrIn_29_TDATA),
    .io_addrIn_30_TREADY(syncSide_io_addrIn_30_TREADY),
    .io_addrIn_30_TVALID(syncSide_io_addrIn_30_TVALID),
    .io_addrIn_30_TDATA(syncSide_io_addrIn_30_TDATA),
    .io_addrIn_31_TREADY(syncSide_io_addrIn_31_TREADY),
    .io_addrIn_31_TVALID(syncSide_io_addrIn_31_TVALID),
    .io_addrIn_31_TDATA(syncSide_io_addrIn_31_TDATA),
    .io_addrIn_32_TREADY(syncSide_io_addrIn_32_TREADY),
    .io_addrIn_32_TVALID(syncSide_io_addrIn_32_TVALID),
    .io_addrIn_32_TDATA(syncSide_io_addrIn_32_TDATA),
    .io_addrIn_33_TREADY(syncSide_io_addrIn_33_TREADY),
    .io_addrIn_33_TVALID(syncSide_io_addrIn_33_TVALID),
    .io_addrIn_33_TDATA(syncSide_io_addrIn_33_TDATA),
    .io_addrIn_34_TREADY(syncSide_io_addrIn_34_TREADY),
    .io_addrIn_34_TVALID(syncSide_io_addrIn_34_TVALID),
    .io_addrIn_34_TDATA(syncSide_io_addrIn_34_TDATA),
    .io_addrIn_35_TREADY(syncSide_io_addrIn_35_TREADY),
    .io_addrIn_35_TVALID(syncSide_io_addrIn_35_TVALID),
    .io_addrIn_35_TDATA(syncSide_io_addrIn_35_TDATA),
    .io_addrIn_36_TREADY(syncSide_io_addrIn_36_TREADY),
    .io_addrIn_36_TVALID(syncSide_io_addrIn_36_TVALID),
    .io_addrIn_36_TDATA(syncSide_io_addrIn_36_TDATA),
    .io_addrIn_37_TREADY(syncSide_io_addrIn_37_TREADY),
    .io_addrIn_37_TVALID(syncSide_io_addrIn_37_TVALID),
    .io_addrIn_37_TDATA(syncSide_io_addrIn_37_TDATA),
    .io_addrIn_38_TREADY(syncSide_io_addrIn_38_TREADY),
    .io_addrIn_38_TVALID(syncSide_io_addrIn_38_TVALID),
    .io_addrIn_38_TDATA(syncSide_io_addrIn_38_TDATA),
    .io_addrIn_39_TREADY(syncSide_io_addrIn_39_TREADY),
    .io_addrIn_39_TVALID(syncSide_io_addrIn_39_TVALID),
    .io_addrIn_39_TDATA(syncSide_io_addrIn_39_TDATA),
    .io_addrIn_40_TREADY(syncSide_io_addrIn_40_TREADY),
    .io_addrIn_40_TVALID(syncSide_io_addrIn_40_TVALID),
    .io_addrIn_40_TDATA(syncSide_io_addrIn_40_TDATA),
    .io_addrIn_41_TREADY(syncSide_io_addrIn_41_TREADY),
    .io_addrIn_41_TVALID(syncSide_io_addrIn_41_TVALID),
    .io_addrIn_41_TDATA(syncSide_io_addrIn_41_TDATA),
    .io_addrIn_42_TREADY(syncSide_io_addrIn_42_TREADY),
    .io_addrIn_42_TVALID(syncSide_io_addrIn_42_TVALID),
    .io_addrIn_42_TDATA(syncSide_io_addrIn_42_TDATA),
    .io_addrIn_43_TREADY(syncSide_io_addrIn_43_TREADY),
    .io_addrIn_43_TVALID(syncSide_io_addrIn_43_TVALID),
    .io_addrIn_43_TDATA(syncSide_io_addrIn_43_TDATA),
    .io_addrIn_44_TREADY(syncSide_io_addrIn_44_TREADY),
    .io_addrIn_44_TVALID(syncSide_io_addrIn_44_TVALID),
    .io_addrIn_44_TDATA(syncSide_io_addrIn_44_TDATA),
    .io_addrIn_45_TREADY(syncSide_io_addrIn_45_TREADY),
    .io_addrIn_45_TVALID(syncSide_io_addrIn_45_TVALID),
    .io_addrIn_45_TDATA(syncSide_io_addrIn_45_TDATA),
    .io_addrIn_46_TREADY(syncSide_io_addrIn_46_TREADY),
    .io_addrIn_46_TVALID(syncSide_io_addrIn_46_TVALID),
    .io_addrIn_46_TDATA(syncSide_io_addrIn_46_TDATA),
    .io_addrIn_47_TREADY(syncSide_io_addrIn_47_TREADY),
    .io_addrIn_47_TVALID(syncSide_io_addrIn_47_TVALID),
    .io_addrIn_47_TDATA(syncSide_io_addrIn_47_TDATA),
    .io_addrIn_48_TREADY(syncSide_io_addrIn_48_TREADY),
    .io_addrIn_48_TVALID(syncSide_io_addrIn_48_TVALID),
    .io_addrIn_48_TDATA(syncSide_io_addrIn_48_TDATA),
    .io_addrIn_49_TREADY(syncSide_io_addrIn_49_TREADY),
    .io_addrIn_49_TVALID(syncSide_io_addrIn_49_TVALID),
    .io_addrIn_49_TDATA(syncSide_io_addrIn_49_TDATA),
    .io_addrIn_50_TREADY(syncSide_io_addrIn_50_TREADY),
    .io_addrIn_50_TVALID(syncSide_io_addrIn_50_TVALID),
    .io_addrIn_50_TDATA(syncSide_io_addrIn_50_TDATA),
    .io_addrIn_51_TREADY(syncSide_io_addrIn_51_TREADY),
    .io_addrIn_51_TVALID(syncSide_io_addrIn_51_TVALID),
    .io_addrIn_51_TDATA(syncSide_io_addrIn_51_TDATA),
    .io_addrIn_52_TREADY(syncSide_io_addrIn_52_TREADY),
    .io_addrIn_52_TVALID(syncSide_io_addrIn_52_TVALID),
    .io_addrIn_52_TDATA(syncSide_io_addrIn_52_TDATA),
    .io_addrIn_53_TREADY(syncSide_io_addrIn_53_TREADY),
    .io_addrIn_53_TVALID(syncSide_io_addrIn_53_TVALID),
    .io_addrIn_53_TDATA(syncSide_io_addrIn_53_TDATA),
    .io_addrIn_54_TREADY(syncSide_io_addrIn_54_TREADY),
    .io_addrIn_54_TVALID(syncSide_io_addrIn_54_TVALID),
    .io_addrIn_54_TDATA(syncSide_io_addrIn_54_TDATA),
    .io_addrIn_55_TREADY(syncSide_io_addrIn_55_TREADY),
    .io_addrIn_55_TVALID(syncSide_io_addrIn_55_TVALID),
    .io_addrIn_55_TDATA(syncSide_io_addrIn_55_TDATA),
    .io_addrIn_56_TREADY(syncSide_io_addrIn_56_TREADY),
    .io_addrIn_56_TVALID(syncSide_io_addrIn_56_TVALID),
    .io_addrIn_56_TDATA(syncSide_io_addrIn_56_TDATA),
    .io_addrIn_57_TREADY(syncSide_io_addrIn_57_TREADY),
    .io_addrIn_57_TVALID(syncSide_io_addrIn_57_TVALID),
    .io_addrIn_57_TDATA(syncSide_io_addrIn_57_TDATA),
    .io_addrIn_58_TREADY(syncSide_io_addrIn_58_TREADY),
    .io_addrIn_58_TVALID(syncSide_io_addrIn_58_TVALID),
    .io_addrIn_58_TDATA(syncSide_io_addrIn_58_TDATA),
    .io_addrIn_59_TREADY(syncSide_io_addrIn_59_TREADY),
    .io_addrIn_59_TVALID(syncSide_io_addrIn_59_TVALID),
    .io_addrIn_59_TDATA(syncSide_io_addrIn_59_TDATA),
    .io_addrIn_60_TREADY(syncSide_io_addrIn_60_TREADY),
    .io_addrIn_60_TVALID(syncSide_io_addrIn_60_TVALID),
    .io_addrIn_60_TDATA(syncSide_io_addrIn_60_TDATA),
    .io_addrIn_61_TREADY(syncSide_io_addrIn_61_TREADY),
    .io_addrIn_61_TVALID(syncSide_io_addrIn_61_TVALID),
    .io_addrIn_61_TDATA(syncSide_io_addrIn_61_TDATA),
    .io_addrIn_62_TREADY(syncSide_io_addrIn_62_TREADY),
    .io_addrIn_62_TVALID(syncSide_io_addrIn_62_TVALID),
    .io_addrIn_62_TDATA(syncSide_io_addrIn_62_TDATA),
    .io_addrIn_63_TREADY(syncSide_io_addrIn_63_TREADY),
    .io_addrIn_63_TVALID(syncSide_io_addrIn_63_TVALID),
    .io_addrIn_63_TDATA(syncSide_io_addrIn_63_TDATA),
    .io_axi_full_argRoute_0_ARREADY(syncSide_io_axi_full_argRoute_0_ARREADY),
    .io_axi_full_argRoute_0_ARVALID(syncSide_io_axi_full_argRoute_0_ARVALID),
    .io_axi_full_argRoute_0_ARADDR(syncSide_io_axi_full_argRoute_0_ARADDR),
    .io_axi_full_argRoute_0_RREADY(syncSide_io_axi_full_argRoute_0_RREADY),
    .io_axi_full_argRoute_0_RVALID(syncSide_io_axi_full_argRoute_0_RVALID),
    .io_axi_full_argRoute_0_RDATA(syncSide_io_axi_full_argRoute_0_RDATA),
    .io_axi_full_argRoute_0_AWREADY(syncSide_io_axi_full_argRoute_0_AWREADY),
    .io_axi_full_argRoute_0_AWVALID(syncSide_io_axi_full_argRoute_0_AWVALID),
    .io_axi_full_argRoute_0_AWADDR(syncSide_io_axi_full_argRoute_0_AWADDR),
    .io_axi_full_argRoute_0_WREADY(syncSide_io_axi_full_argRoute_0_WREADY),
    .io_axi_full_argRoute_0_WVALID(syncSide_io_axi_full_argRoute_0_WVALID),
    .io_axi_full_argRoute_0_WDATA(syncSide_io_axi_full_argRoute_0_WDATA),
    .io_axi_full_argRoute_0_BVALID(syncSide_io_axi_full_argRoute_0_BVALID),
    .io_axi_full_argRoute_1_ARREADY(syncSide_io_axi_full_argRoute_1_ARREADY),
    .io_axi_full_argRoute_1_ARVALID(syncSide_io_axi_full_argRoute_1_ARVALID),
    .io_axi_full_argRoute_1_ARADDR(syncSide_io_axi_full_argRoute_1_ARADDR),
    .io_axi_full_argRoute_1_RREADY(syncSide_io_axi_full_argRoute_1_RREADY),
    .io_axi_full_argRoute_1_RVALID(syncSide_io_axi_full_argRoute_1_RVALID),
    .io_axi_full_argRoute_1_RDATA(syncSide_io_axi_full_argRoute_1_RDATA),
    .io_axi_full_argRoute_1_AWREADY(syncSide_io_axi_full_argRoute_1_AWREADY),
    .io_axi_full_argRoute_1_AWVALID(syncSide_io_axi_full_argRoute_1_AWVALID),
    .io_axi_full_argRoute_1_AWADDR(syncSide_io_axi_full_argRoute_1_AWADDR),
    .io_axi_full_argRoute_1_WREADY(syncSide_io_axi_full_argRoute_1_WREADY),
    .io_axi_full_argRoute_1_WVALID(syncSide_io_axi_full_argRoute_1_WVALID),
    .io_axi_full_argRoute_1_WDATA(syncSide_io_axi_full_argRoute_1_WDATA),
    .io_axi_full_argRoute_1_BVALID(syncSide_io_axi_full_argRoute_1_BVALID),
    .io_axi_full_argRoute_2_ARREADY(syncSide_io_axi_full_argRoute_2_ARREADY),
    .io_axi_full_argRoute_2_ARVALID(syncSide_io_axi_full_argRoute_2_ARVALID),
    .io_axi_full_argRoute_2_ARADDR(syncSide_io_axi_full_argRoute_2_ARADDR),
    .io_axi_full_argRoute_2_RREADY(syncSide_io_axi_full_argRoute_2_RREADY),
    .io_axi_full_argRoute_2_RVALID(syncSide_io_axi_full_argRoute_2_RVALID),
    .io_axi_full_argRoute_2_RDATA(syncSide_io_axi_full_argRoute_2_RDATA),
    .io_axi_full_argRoute_3_ARREADY(syncSide_io_axi_full_argRoute_3_ARREADY),
    .io_axi_full_argRoute_3_ARVALID(syncSide_io_axi_full_argRoute_3_ARVALID),
    .io_axi_full_argRoute_3_ARADDR(syncSide_io_axi_full_argRoute_3_ARADDR),
    .io_axi_full_argRoute_3_RREADY(syncSide_io_axi_full_argRoute_3_RREADY),
    .io_axi_full_argRoute_3_RVALID(syncSide_io_axi_full_argRoute_3_RVALID),
    .io_axi_full_argRoute_3_RDATA(syncSide_io_axi_full_argRoute_3_RDATA),
    .connStealNtw_0_ctrl_serveStealReq_ready(syncSide_connStealNtw_0_ctrl_serveStealReq_ready),
    .connStealNtw_0_ctrl_serveStealReq_valid(syncSide_connStealNtw_0_ctrl_serveStealReq_valid),
    .connStealNtw_0_data_qOutTask_ready(syncSide_connStealNtw_0_data_qOutTask_ready),
    .connStealNtw_0_data_qOutTask_valid(syncSide_connStealNtw_0_data_qOutTask_valid),
    .connStealNtw_0_data_qOutTask_bits(syncSide_connStealNtw_0_data_qOutTask_bits),
    .connStealNtw_1_ctrl_serveStealReq_ready(syncSide_connStealNtw_1_ctrl_serveStealReq_ready),
    .connStealNtw_1_ctrl_serveStealReq_valid(syncSide_connStealNtw_1_ctrl_serveStealReq_valid),
    .connStealNtw_1_data_qOutTask_ready(syncSide_connStealNtw_1_data_qOutTask_ready),
    .connStealNtw_1_data_qOutTask_valid(syncSide_connStealNtw_1_data_qOutTask_valid),
    .connStealNtw_1_data_qOutTask_bits(syncSide_connStealNtw_1_data_qOutTask_bits)
  );
  assign task_stealSide_axi_mgmt_vss_0_ARREADY = stealSide_io_axi_mgmt_vss_0_ARREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_axi_mgmt_vss_0_RVALID = stealSide_io_axi_mgmt_vss_0_RVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_axi_mgmt_vss_0_RDATA = stealSide_io_axi_mgmt_vss_0_RDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_axi_mgmt_vss_0_RRESP = 2'h0; // @[fullSysGen.scala 246:23]
  assign task_stealSide_axi_mgmt_vss_0_AWREADY = stealSide_io_axi_mgmt_vss_0_AWREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_axi_mgmt_vss_0_WREADY = stealSide_io_axi_mgmt_vss_0_WREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_axi_mgmt_vss_0_BVALID = stealSide_io_axi_mgmt_vss_0_BVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_axi_mgmt_vss_0_BRESP = 2'h0; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_ARVALID = stealSide_io_vss_axi_full_0_ARVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_ARID = 4'h0; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_ARADDR = stealSide_io_vss_axi_full_0_ARADDR; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_ARLEN = stealSide_io_vss_axi_full_0_ARLEN; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_ARSIZE = 3'h5; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_ARBURST = 2'h1; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_ARLOCK = 1'h0; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_ARCACHE = 4'h0; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_ARPROT = 3'h0; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_ARQOS = 4'h0; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_ARREGION = 4'h0; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_RREADY = stealSide_io_vss_axi_full_0_RREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_AWVALID = stealSide_io_vss_axi_full_0_AWVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_AWID = 4'h0; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_AWADDR = stealSide_io_vss_axi_full_0_AWADDR; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_AWLEN = stealSide_io_vss_axi_full_0_AWLEN; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_AWSIZE = 3'h5; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_AWBURST = 2'h1; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_AWLOCK = 1'h0; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_AWCACHE = 4'h0; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_AWPROT = 3'h0; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_AWQOS = 4'h0; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_AWREGION = 4'h0; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_WVALID = stealSide_io_vss_axi_full_0_WVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_WID = 4'h0; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_WDATA = stealSide_io_vss_axi_full_0_WDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_WSTRB = 32'hffffffff; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_WLAST = stealSide_io_vss_axi_full_0_WLAST; // @[fullSysGen.scala 246:23]
  assign task_stealSide_vss_axi_full_0_BREADY = 1'h1; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_0_TVALID = stealSide_io_taskOut_0_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_0_TDATA = stealSide_io_taskOut_0_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_1_TVALID = stealSide_io_taskOut_1_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_1_TDATA = stealSide_io_taskOut_1_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_2_TVALID = stealSide_io_taskOut_2_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_2_TDATA = stealSide_io_taskOut_2_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_3_TVALID = stealSide_io_taskOut_3_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_3_TDATA = stealSide_io_taskOut_3_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_4_TVALID = stealSide_io_taskOut_4_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_4_TDATA = stealSide_io_taskOut_4_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_5_TVALID = stealSide_io_taskOut_5_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_5_TDATA = stealSide_io_taskOut_5_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_6_TVALID = stealSide_io_taskOut_6_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_6_TDATA = stealSide_io_taskOut_6_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_7_TVALID = stealSide_io_taskOut_7_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_7_TDATA = stealSide_io_taskOut_7_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_8_TVALID = stealSide_io_taskOut_8_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_8_TDATA = stealSide_io_taskOut_8_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_9_TVALID = stealSide_io_taskOut_9_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_9_TDATA = stealSide_io_taskOut_9_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_10_TVALID = stealSide_io_taskOut_10_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_10_TDATA = stealSide_io_taskOut_10_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_11_TVALID = stealSide_io_taskOut_11_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_11_TDATA = stealSide_io_taskOut_11_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_12_TVALID = stealSide_io_taskOut_12_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_12_TDATA = stealSide_io_taskOut_12_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_13_TVALID = stealSide_io_taskOut_13_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_13_TDATA = stealSide_io_taskOut_13_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_14_TVALID = stealSide_io_taskOut_14_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_14_TDATA = stealSide_io_taskOut_14_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_15_TVALID = stealSide_io_taskOut_15_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_15_TDATA = stealSide_io_taskOut_15_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_16_TVALID = stealSide_io_taskOut_16_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_16_TDATA = stealSide_io_taskOut_16_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_17_TVALID = stealSide_io_taskOut_17_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_17_TDATA = stealSide_io_taskOut_17_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_18_TVALID = stealSide_io_taskOut_18_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_18_TDATA = stealSide_io_taskOut_18_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_19_TVALID = stealSide_io_taskOut_19_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_19_TDATA = stealSide_io_taskOut_19_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_20_TVALID = stealSide_io_taskOut_20_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_20_TDATA = stealSide_io_taskOut_20_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_21_TVALID = stealSide_io_taskOut_21_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_21_TDATA = stealSide_io_taskOut_21_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_22_TVALID = stealSide_io_taskOut_22_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_22_TDATA = stealSide_io_taskOut_22_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_23_TVALID = stealSide_io_taskOut_23_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_23_TDATA = stealSide_io_taskOut_23_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_24_TVALID = stealSide_io_taskOut_24_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_24_TDATA = stealSide_io_taskOut_24_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_25_TVALID = stealSide_io_taskOut_25_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_25_TDATA = stealSide_io_taskOut_25_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_26_TVALID = stealSide_io_taskOut_26_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_26_TDATA = stealSide_io_taskOut_26_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_27_TVALID = stealSide_io_taskOut_27_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_27_TDATA = stealSide_io_taskOut_27_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_28_TVALID = stealSide_io_taskOut_28_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_28_TDATA = stealSide_io_taskOut_28_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_29_TVALID = stealSide_io_taskOut_29_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_29_TDATA = stealSide_io_taskOut_29_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_30_TVALID = stealSide_io_taskOut_30_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_30_TDATA = stealSide_io_taskOut_30_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_31_TVALID = stealSide_io_taskOut_31_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_31_TDATA = stealSide_io_taskOut_31_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_32_TVALID = stealSide_io_taskOut_32_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_32_TDATA = stealSide_io_taskOut_32_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_33_TVALID = stealSide_io_taskOut_33_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_33_TDATA = stealSide_io_taskOut_33_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_34_TVALID = stealSide_io_taskOut_34_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_34_TDATA = stealSide_io_taskOut_34_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_35_TVALID = stealSide_io_taskOut_35_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_35_TDATA = stealSide_io_taskOut_35_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_36_TVALID = stealSide_io_taskOut_36_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_36_TDATA = stealSide_io_taskOut_36_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_37_TVALID = stealSide_io_taskOut_37_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_37_TDATA = stealSide_io_taskOut_37_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_38_TVALID = stealSide_io_taskOut_38_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_38_TDATA = stealSide_io_taskOut_38_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_39_TVALID = stealSide_io_taskOut_39_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_39_TDATA = stealSide_io_taskOut_39_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_40_TVALID = stealSide_io_taskOut_40_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_40_TDATA = stealSide_io_taskOut_40_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_41_TVALID = stealSide_io_taskOut_41_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_41_TDATA = stealSide_io_taskOut_41_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_42_TVALID = stealSide_io_taskOut_42_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_42_TDATA = stealSide_io_taskOut_42_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_43_TVALID = stealSide_io_taskOut_43_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_43_TDATA = stealSide_io_taskOut_43_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_44_TVALID = stealSide_io_taskOut_44_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_44_TDATA = stealSide_io_taskOut_44_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_45_TVALID = stealSide_io_taskOut_45_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_45_TDATA = stealSide_io_taskOut_45_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_46_TVALID = stealSide_io_taskOut_46_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_46_TDATA = stealSide_io_taskOut_46_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_47_TVALID = stealSide_io_taskOut_47_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_47_TDATA = stealSide_io_taskOut_47_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_48_TVALID = stealSide_io_taskOut_48_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_48_TDATA = stealSide_io_taskOut_48_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_49_TVALID = stealSide_io_taskOut_49_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_49_TDATA = stealSide_io_taskOut_49_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_50_TVALID = stealSide_io_taskOut_50_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_50_TDATA = stealSide_io_taskOut_50_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_51_TVALID = stealSide_io_taskOut_51_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_51_TDATA = stealSide_io_taskOut_51_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_52_TVALID = stealSide_io_taskOut_52_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_52_TDATA = stealSide_io_taskOut_52_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_53_TVALID = stealSide_io_taskOut_53_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_53_TDATA = stealSide_io_taskOut_53_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_54_TVALID = stealSide_io_taskOut_54_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_54_TDATA = stealSide_io_taskOut_54_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_55_TVALID = stealSide_io_taskOut_55_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_55_TDATA = stealSide_io_taskOut_55_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_56_TVALID = stealSide_io_taskOut_56_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_56_TDATA = stealSide_io_taskOut_56_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_57_TVALID = stealSide_io_taskOut_57_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_57_TDATA = stealSide_io_taskOut_57_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_58_TVALID = stealSide_io_taskOut_58_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_58_TDATA = stealSide_io_taskOut_58_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_59_TVALID = stealSide_io_taskOut_59_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_59_TDATA = stealSide_io_taskOut_59_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_60_TVALID = stealSide_io_taskOut_60_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_60_TDATA = stealSide_io_taskOut_60_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_61_TVALID = stealSide_io_taskOut_61_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_61_TDATA = stealSide_io_taskOut_61_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_62_TVALID = stealSide_io_taskOut_62_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_62_TDATA = stealSide_io_taskOut_62_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_63_TVALID = stealSide_io_taskOut_63_TVALID; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskOut_63_TDATA = stealSide_io_taskOut_63_TDATA; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_0_TREADY = stealSide_io_taskIn_0_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_1_TREADY = stealSide_io_taskIn_1_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_2_TREADY = stealSide_io_taskIn_2_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_3_TREADY = stealSide_io_taskIn_3_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_4_TREADY = stealSide_io_taskIn_4_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_5_TREADY = stealSide_io_taskIn_5_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_6_TREADY = stealSide_io_taskIn_6_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_7_TREADY = stealSide_io_taskIn_7_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_8_TREADY = stealSide_io_taskIn_8_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_9_TREADY = stealSide_io_taskIn_9_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_10_TREADY = stealSide_io_taskIn_10_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_11_TREADY = stealSide_io_taskIn_11_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_12_TREADY = stealSide_io_taskIn_12_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_13_TREADY = stealSide_io_taskIn_13_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_14_TREADY = stealSide_io_taskIn_14_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_15_TREADY = stealSide_io_taskIn_15_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_16_TREADY = stealSide_io_taskIn_16_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_17_TREADY = stealSide_io_taskIn_17_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_18_TREADY = stealSide_io_taskIn_18_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_19_TREADY = stealSide_io_taskIn_19_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_20_TREADY = stealSide_io_taskIn_20_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_21_TREADY = stealSide_io_taskIn_21_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_22_TREADY = stealSide_io_taskIn_22_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_23_TREADY = stealSide_io_taskIn_23_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_24_TREADY = stealSide_io_taskIn_24_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_25_TREADY = stealSide_io_taskIn_25_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_26_TREADY = stealSide_io_taskIn_26_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_27_TREADY = stealSide_io_taskIn_27_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_28_TREADY = stealSide_io_taskIn_28_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_29_TREADY = stealSide_io_taskIn_29_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_30_TREADY = stealSide_io_taskIn_30_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_31_TREADY = stealSide_io_taskIn_31_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_32_TREADY = stealSide_io_taskIn_32_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_33_TREADY = stealSide_io_taskIn_33_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_34_TREADY = stealSide_io_taskIn_34_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_35_TREADY = stealSide_io_taskIn_35_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_36_TREADY = stealSide_io_taskIn_36_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_37_TREADY = stealSide_io_taskIn_37_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_38_TREADY = stealSide_io_taskIn_38_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_39_TREADY = stealSide_io_taskIn_39_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_40_TREADY = stealSide_io_taskIn_40_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_41_TREADY = stealSide_io_taskIn_41_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_42_TREADY = stealSide_io_taskIn_42_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_43_TREADY = stealSide_io_taskIn_43_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_44_TREADY = stealSide_io_taskIn_44_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_45_TREADY = stealSide_io_taskIn_45_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_46_TREADY = stealSide_io_taskIn_46_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_47_TREADY = stealSide_io_taskIn_47_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_48_TREADY = stealSide_io_taskIn_48_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_49_TREADY = stealSide_io_taskIn_49_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_50_TREADY = stealSide_io_taskIn_50_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_51_TREADY = stealSide_io_taskIn_51_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_52_TREADY = stealSide_io_taskIn_52_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_53_TREADY = stealSide_io_taskIn_53_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_54_TREADY = stealSide_io_taskIn_54_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_55_TREADY = stealSide_io_taskIn_55_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_56_TREADY = stealSide_io_taskIn_56_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_57_TREADY = stealSide_io_taskIn_57_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_58_TREADY = stealSide_io_taskIn_58_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_59_TREADY = stealSide_io_taskIn_59_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_60_TREADY = stealSide_io_taskIn_60_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_61_TREADY = stealSide_io_taskIn_61_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_62_TREADY = stealSide_io_taskIn_62_TREADY; // @[fullSysGen.scala 246:23]
  assign task_stealSide_taskIn_63_TREADY = stealSide_io_taskIn_63_TREADY; // @[fullSysGen.scala 246:23]
  assign task_continuationAllocationSide_contOut_0_TVALID = continuationAllocationSide_io_contOut_0_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_0_TDATA = continuationAllocationSide_io_contOut_0_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_1_TVALID = continuationAllocationSide_io_contOut_1_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_1_TDATA = continuationAllocationSide_io_contOut_1_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_2_TVALID = continuationAllocationSide_io_contOut_2_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_2_TDATA = continuationAllocationSide_io_contOut_2_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_3_TVALID = continuationAllocationSide_io_contOut_3_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_3_TDATA = continuationAllocationSide_io_contOut_3_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_4_TVALID = continuationAllocationSide_io_contOut_4_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_4_TDATA = continuationAllocationSide_io_contOut_4_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_5_TVALID = continuationAllocationSide_io_contOut_5_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_5_TDATA = continuationAllocationSide_io_contOut_5_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_6_TVALID = continuationAllocationSide_io_contOut_6_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_6_TDATA = continuationAllocationSide_io_contOut_6_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_7_TVALID = continuationAllocationSide_io_contOut_7_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_7_TDATA = continuationAllocationSide_io_contOut_7_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_8_TVALID = continuationAllocationSide_io_contOut_8_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_8_TDATA = continuationAllocationSide_io_contOut_8_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_9_TVALID = continuationAllocationSide_io_contOut_9_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_9_TDATA = continuationAllocationSide_io_contOut_9_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_10_TVALID = continuationAllocationSide_io_contOut_10_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_10_TDATA = continuationAllocationSide_io_contOut_10_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_11_TVALID = continuationAllocationSide_io_contOut_11_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_11_TDATA = continuationAllocationSide_io_contOut_11_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_12_TVALID = continuationAllocationSide_io_contOut_12_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_12_TDATA = continuationAllocationSide_io_contOut_12_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_13_TVALID = continuationAllocationSide_io_contOut_13_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_13_TDATA = continuationAllocationSide_io_contOut_13_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_14_TVALID = continuationAllocationSide_io_contOut_14_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_14_TDATA = continuationAllocationSide_io_contOut_14_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_15_TVALID = continuationAllocationSide_io_contOut_15_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_15_TDATA = continuationAllocationSide_io_contOut_15_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_16_TVALID = continuationAllocationSide_io_contOut_16_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_16_TDATA = continuationAllocationSide_io_contOut_16_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_17_TVALID = continuationAllocationSide_io_contOut_17_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_17_TDATA = continuationAllocationSide_io_contOut_17_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_18_TVALID = continuationAllocationSide_io_contOut_18_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_18_TDATA = continuationAllocationSide_io_contOut_18_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_19_TVALID = continuationAllocationSide_io_contOut_19_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_19_TDATA = continuationAllocationSide_io_contOut_19_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_20_TVALID = continuationAllocationSide_io_contOut_20_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_20_TDATA = continuationAllocationSide_io_contOut_20_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_21_TVALID = continuationAllocationSide_io_contOut_21_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_21_TDATA = continuationAllocationSide_io_contOut_21_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_22_TVALID = continuationAllocationSide_io_contOut_22_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_22_TDATA = continuationAllocationSide_io_contOut_22_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_23_TVALID = continuationAllocationSide_io_contOut_23_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_23_TDATA = continuationAllocationSide_io_contOut_23_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_24_TVALID = continuationAllocationSide_io_contOut_24_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_24_TDATA = continuationAllocationSide_io_contOut_24_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_25_TVALID = continuationAllocationSide_io_contOut_25_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_25_TDATA = continuationAllocationSide_io_contOut_25_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_26_TVALID = continuationAllocationSide_io_contOut_26_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_26_TDATA = continuationAllocationSide_io_contOut_26_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_27_TVALID = continuationAllocationSide_io_contOut_27_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_27_TDATA = continuationAllocationSide_io_contOut_27_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_28_TVALID = continuationAllocationSide_io_contOut_28_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_28_TDATA = continuationAllocationSide_io_contOut_28_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_29_TVALID = continuationAllocationSide_io_contOut_29_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_29_TDATA = continuationAllocationSide_io_contOut_29_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_30_TVALID = continuationAllocationSide_io_contOut_30_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_30_TDATA = continuationAllocationSide_io_contOut_30_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_31_TVALID = continuationAllocationSide_io_contOut_31_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_31_TDATA = continuationAllocationSide_io_contOut_31_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_32_TVALID = continuationAllocationSide_io_contOut_32_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_32_TDATA = continuationAllocationSide_io_contOut_32_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_33_TVALID = continuationAllocationSide_io_contOut_33_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_33_TDATA = continuationAllocationSide_io_contOut_33_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_34_TVALID = continuationAllocationSide_io_contOut_34_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_34_TDATA = continuationAllocationSide_io_contOut_34_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_35_TVALID = continuationAllocationSide_io_contOut_35_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_35_TDATA = continuationAllocationSide_io_contOut_35_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_36_TVALID = continuationAllocationSide_io_contOut_36_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_36_TDATA = continuationAllocationSide_io_contOut_36_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_37_TVALID = continuationAllocationSide_io_contOut_37_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_37_TDATA = continuationAllocationSide_io_contOut_37_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_38_TVALID = continuationAllocationSide_io_contOut_38_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_38_TDATA = continuationAllocationSide_io_contOut_38_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_39_TVALID = continuationAllocationSide_io_contOut_39_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_39_TDATA = continuationAllocationSide_io_contOut_39_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_40_TVALID = continuationAllocationSide_io_contOut_40_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_40_TDATA = continuationAllocationSide_io_contOut_40_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_41_TVALID = continuationAllocationSide_io_contOut_41_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_41_TDATA = continuationAllocationSide_io_contOut_41_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_42_TVALID = continuationAllocationSide_io_contOut_42_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_42_TDATA = continuationAllocationSide_io_contOut_42_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_43_TVALID = continuationAllocationSide_io_contOut_43_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_43_TDATA = continuationAllocationSide_io_contOut_43_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_44_TVALID = continuationAllocationSide_io_contOut_44_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_44_TDATA = continuationAllocationSide_io_contOut_44_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_45_TVALID = continuationAllocationSide_io_contOut_45_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_45_TDATA = continuationAllocationSide_io_contOut_45_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_46_TVALID = continuationAllocationSide_io_contOut_46_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_46_TDATA = continuationAllocationSide_io_contOut_46_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_47_TVALID = continuationAllocationSide_io_contOut_47_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_47_TDATA = continuationAllocationSide_io_contOut_47_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_48_TVALID = continuationAllocationSide_io_contOut_48_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_48_TDATA = continuationAllocationSide_io_contOut_48_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_49_TVALID = continuationAllocationSide_io_contOut_49_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_49_TDATA = continuationAllocationSide_io_contOut_49_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_50_TVALID = continuationAllocationSide_io_contOut_50_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_50_TDATA = continuationAllocationSide_io_contOut_50_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_51_TVALID = continuationAllocationSide_io_contOut_51_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_51_TDATA = continuationAllocationSide_io_contOut_51_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_52_TVALID = continuationAllocationSide_io_contOut_52_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_52_TDATA = continuationAllocationSide_io_contOut_52_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_53_TVALID = continuationAllocationSide_io_contOut_53_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_53_TDATA = continuationAllocationSide_io_contOut_53_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_54_TVALID = continuationAllocationSide_io_contOut_54_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_54_TDATA = continuationAllocationSide_io_contOut_54_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_55_TVALID = continuationAllocationSide_io_contOut_55_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_55_TDATA = continuationAllocationSide_io_contOut_55_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_56_TVALID = continuationAllocationSide_io_contOut_56_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_56_TDATA = continuationAllocationSide_io_contOut_56_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_57_TVALID = continuationAllocationSide_io_contOut_57_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_57_TDATA = continuationAllocationSide_io_contOut_57_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_58_TVALID = continuationAllocationSide_io_contOut_58_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_58_TDATA = continuationAllocationSide_io_contOut_58_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_59_TVALID = continuationAllocationSide_io_contOut_59_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_59_TDATA = continuationAllocationSide_io_contOut_59_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_60_TVALID = continuationAllocationSide_io_contOut_60_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_60_TDATA = continuationAllocationSide_io_contOut_60_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_61_TVALID = continuationAllocationSide_io_contOut_61_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_61_TDATA = continuationAllocationSide_io_contOut_61_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_62_TVALID = continuationAllocationSide_io_contOut_62_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_62_TDATA = continuationAllocationSide_io_contOut_62_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_63_TVALID = continuationAllocationSide_io_contOut_63_TVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_contOut_63_TDATA = continuationAllocationSide_io_contOut_63_TDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_axi_mgmt_vcas_0_ARREADY = continuationAllocationSide_io_axi_mgmt_vcas_0_ARREADY
    ; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_axi_mgmt_vcas_0_RVALID = continuationAllocationSide_io_axi_mgmt_vcas_0_RVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_axi_mgmt_vcas_0_RDATA = continuationAllocationSide_io_axi_mgmt_vcas_0_RDATA; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_axi_mgmt_vcas_0_RRESP = 2'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_axi_mgmt_vcas_0_AWREADY = continuationAllocationSide_io_axi_mgmt_vcas_0_AWREADY
    ; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_axi_mgmt_vcas_0_WREADY = continuationAllocationSide_io_axi_mgmt_vcas_0_WREADY; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_axi_mgmt_vcas_0_BVALID = continuationAllocationSide_io_axi_mgmt_vcas_0_BVALID; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_axi_mgmt_vcas_0_BRESP = 2'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_ARVALID = continuationAllocationSide_io_vcas_axi_full_0_ARVALID
    ; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_ARID = 4'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_ARADDR = continuationAllocationSide_io_vcas_axi_full_0_ARADDR; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_ARLEN = 8'hf; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_ARSIZE = 3'h3; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_ARBURST = 2'h1; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_ARLOCK = 1'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_ARCACHE = 4'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_ARPROT = 3'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_ARQOS = 4'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_ARREGION = 4'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_RREADY = continuationAllocationSide_io_vcas_axi_full_0_RREADY; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_AWVALID = 1'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_AWID = 4'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_AWADDR = 64'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_AWLEN = 8'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_AWSIZE = 3'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_AWBURST = 2'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_AWLOCK = 1'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_AWCACHE = 4'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_AWPROT = 3'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_AWQOS = 4'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_AWREGION = 4'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_WVALID = 1'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_WID = 4'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_WDATA = 64'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_WSTRB = 8'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_WLAST = 1'h0; // @[fullSysGen.scala 282:42]
  assign task_continuationAllocationSide_vcas_axi_full_0_BREADY = 1'h0; // @[fullSysGen.scala 282:42]
  assign task_syncSide_addrIn_0_TREADY = syncSide_io_addrIn_0_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_1_TREADY = syncSide_io_addrIn_1_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_2_TREADY = syncSide_io_addrIn_2_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_3_TREADY = syncSide_io_addrIn_3_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_4_TREADY = syncSide_io_addrIn_4_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_5_TREADY = syncSide_io_addrIn_5_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_6_TREADY = syncSide_io_addrIn_6_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_7_TREADY = syncSide_io_addrIn_7_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_8_TREADY = syncSide_io_addrIn_8_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_9_TREADY = syncSide_io_addrIn_9_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_10_TREADY = syncSide_io_addrIn_10_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_11_TREADY = syncSide_io_addrIn_11_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_12_TREADY = syncSide_io_addrIn_12_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_13_TREADY = syncSide_io_addrIn_13_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_14_TREADY = syncSide_io_addrIn_14_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_15_TREADY = syncSide_io_addrIn_15_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_16_TREADY = syncSide_io_addrIn_16_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_17_TREADY = syncSide_io_addrIn_17_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_18_TREADY = syncSide_io_addrIn_18_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_19_TREADY = syncSide_io_addrIn_19_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_20_TREADY = syncSide_io_addrIn_20_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_21_TREADY = syncSide_io_addrIn_21_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_22_TREADY = syncSide_io_addrIn_22_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_23_TREADY = syncSide_io_addrIn_23_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_24_TREADY = syncSide_io_addrIn_24_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_25_TREADY = syncSide_io_addrIn_25_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_26_TREADY = syncSide_io_addrIn_26_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_27_TREADY = syncSide_io_addrIn_27_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_28_TREADY = syncSide_io_addrIn_28_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_29_TREADY = syncSide_io_addrIn_29_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_30_TREADY = syncSide_io_addrIn_30_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_31_TREADY = syncSide_io_addrIn_31_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_32_TREADY = syncSide_io_addrIn_32_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_33_TREADY = syncSide_io_addrIn_33_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_34_TREADY = syncSide_io_addrIn_34_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_35_TREADY = syncSide_io_addrIn_35_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_36_TREADY = syncSide_io_addrIn_36_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_37_TREADY = syncSide_io_addrIn_37_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_38_TREADY = syncSide_io_addrIn_38_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_39_TREADY = syncSide_io_addrIn_39_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_40_TREADY = syncSide_io_addrIn_40_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_41_TREADY = syncSide_io_addrIn_41_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_42_TREADY = syncSide_io_addrIn_42_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_43_TREADY = syncSide_io_addrIn_43_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_44_TREADY = syncSide_io_addrIn_44_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_45_TREADY = syncSide_io_addrIn_45_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_46_TREADY = syncSide_io_addrIn_46_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_47_TREADY = syncSide_io_addrIn_47_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_48_TREADY = syncSide_io_addrIn_48_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_49_TREADY = syncSide_io_addrIn_49_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_50_TREADY = syncSide_io_addrIn_50_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_51_TREADY = syncSide_io_addrIn_51_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_52_TREADY = syncSide_io_addrIn_52_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_53_TREADY = syncSide_io_addrIn_53_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_54_TREADY = syncSide_io_addrIn_54_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_55_TREADY = syncSide_io_addrIn_55_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_56_TREADY = syncSide_io_addrIn_56_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_57_TREADY = syncSide_io_addrIn_57_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_58_TREADY = syncSide_io_addrIn_58_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_59_TREADY = syncSide_io_addrIn_59_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_60_TREADY = syncSide_io_addrIn_60_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_61_TREADY = syncSide_io_addrIn_61_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_62_TREADY = syncSide_io_addrIn_62_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_addrIn_63_TREADY = syncSide_io_addrIn_63_TREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_ARVALID = syncSide_io_axi_full_argRoute_0_ARVALID; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_ARID = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_ARADDR = syncSide_io_axi_full_argRoute_0_ARADDR; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_ARLEN = 8'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_ARSIZE = 3'h2; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_ARBURST = 2'h1; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_ARLOCK = 1'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_ARCACHE = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_ARPROT = 3'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_ARQOS = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_ARREGION = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_RREADY = syncSide_io_axi_full_argRoute_0_RREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_AWVALID = syncSide_io_axi_full_argRoute_0_AWVALID; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_AWID = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_AWADDR = syncSide_io_axi_full_argRoute_0_AWADDR; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_AWLEN = 8'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_AWSIZE = 3'h2; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_AWBURST = 2'h1; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_AWLOCK = 1'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_AWCACHE = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_AWPROT = 3'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_AWQOS = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_AWREGION = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_WVALID = syncSide_io_axi_full_argRoute_0_WVALID; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_WID = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_WDATA = syncSide_io_axi_full_argRoute_0_WDATA; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_WSTRB = 4'hf; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_WLAST = 1'h1; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_0_BREADY = 1'h1; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_ARVALID = syncSide_io_axi_full_argRoute_1_ARVALID; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_ARID = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_ARADDR = syncSide_io_axi_full_argRoute_1_ARADDR; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_ARLEN = 8'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_ARSIZE = 3'h2; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_ARBURST = 2'h1; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_ARLOCK = 1'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_ARCACHE = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_ARPROT = 3'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_ARQOS = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_ARREGION = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_RREADY = syncSide_io_axi_full_argRoute_1_RREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_AWVALID = syncSide_io_axi_full_argRoute_1_AWVALID; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_AWID = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_AWADDR = syncSide_io_axi_full_argRoute_1_AWADDR; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_AWLEN = 8'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_AWSIZE = 3'h2; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_AWBURST = 2'h1; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_AWLOCK = 1'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_AWCACHE = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_AWPROT = 3'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_AWQOS = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_AWREGION = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_WVALID = syncSide_io_axi_full_argRoute_1_WVALID; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_WID = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_WDATA = syncSide_io_axi_full_argRoute_1_WDATA; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_WSTRB = 4'hf; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_WLAST = 1'h1; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_1_BREADY = 1'h1; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_ARVALID = syncSide_io_axi_full_argRoute_2_ARVALID; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_ARID = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_ARADDR = syncSide_io_axi_full_argRoute_2_ARADDR; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_ARLEN = 8'h6; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_ARSIZE = 3'h2; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_ARBURST = 2'h1; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_ARLOCK = 1'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_ARCACHE = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_ARPROT = 3'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_ARQOS = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_ARREGION = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_RREADY = syncSide_io_axi_full_argRoute_2_RREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_AWVALID = 1'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_AWID = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_AWADDR = 64'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_AWLEN = 8'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_AWSIZE = 3'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_AWBURST = 2'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_AWLOCK = 1'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_AWCACHE = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_AWPROT = 3'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_AWQOS = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_AWREGION = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_WVALID = 1'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_WID = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_WDATA = 32'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_WSTRB = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_WLAST = 1'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_2_BREADY = 1'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_ARVALID = syncSide_io_axi_full_argRoute_3_ARVALID; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_ARID = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_ARADDR = syncSide_io_axi_full_argRoute_3_ARADDR; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_ARLEN = 8'h6; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_ARSIZE = 3'h2; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_ARBURST = 2'h1; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_ARLOCK = 1'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_ARCACHE = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_ARPROT = 3'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_ARQOS = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_ARREGION = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_RREADY = syncSide_io_axi_full_argRoute_3_RREADY; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_AWVALID = 1'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_AWID = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_AWADDR = 64'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_AWLEN = 8'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_AWSIZE = 3'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_AWBURST = 2'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_AWLOCK = 1'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_AWCACHE = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_AWPROT = 3'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_AWQOS = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_AWREGION = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_WVALID = 1'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_WID = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_WDATA = 32'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_WSTRB = 4'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_WLAST = 1'h0; // @[fullSysGen.scala 298:24]
  assign task_syncSide_axi_full_argRoute_3_BREADY = 1'h0; // @[fullSysGen.scala 298:24]
  assign stealSide_clock = clock;
  assign stealSide_reset = reset;
  assign stealSide_io_axi_mgmt_vss_0_ARVALID = task_stealSide_axi_mgmt_vss_0_ARVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_axi_mgmt_vss_0_ARADDR = task_stealSide_axi_mgmt_vss_0_ARADDR; // @[fullSysGen.scala 246:23]
  assign stealSide_io_axi_mgmt_vss_0_RREADY = task_stealSide_axi_mgmt_vss_0_RREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_axi_mgmt_vss_0_AWVALID = task_stealSide_axi_mgmt_vss_0_AWVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_axi_mgmt_vss_0_AWADDR = task_stealSide_axi_mgmt_vss_0_AWADDR; // @[fullSysGen.scala 246:23]
  assign stealSide_io_axi_mgmt_vss_0_WVALID = task_stealSide_axi_mgmt_vss_0_WVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_axi_mgmt_vss_0_WDATA = task_stealSide_axi_mgmt_vss_0_WDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_axi_mgmt_vss_0_WSTRB = task_stealSide_axi_mgmt_vss_0_WSTRB; // @[fullSysGen.scala 246:23]
  assign stealSide_io_axi_mgmt_vss_0_BREADY = task_stealSide_axi_mgmt_vss_0_BREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_vss_axi_full_0_ARREADY = task_stealSide_vss_axi_full_0_ARREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_vss_axi_full_0_RVALID = task_stealSide_vss_axi_full_0_RVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_vss_axi_full_0_RDATA = task_stealSide_vss_axi_full_0_RDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_vss_axi_full_0_AWREADY = task_stealSide_vss_axi_full_0_AWREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_vss_axi_full_0_WREADY = task_stealSide_vss_axi_full_0_WREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_vss_axi_full_0_BVALID = task_stealSide_vss_axi_full_0_BVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_0_TREADY = task_stealSide_taskOut_0_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_1_TREADY = task_stealSide_taskOut_1_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_2_TREADY = task_stealSide_taskOut_2_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_3_TREADY = task_stealSide_taskOut_3_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_4_TREADY = task_stealSide_taskOut_4_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_5_TREADY = task_stealSide_taskOut_5_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_6_TREADY = task_stealSide_taskOut_6_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_7_TREADY = task_stealSide_taskOut_7_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_8_TREADY = task_stealSide_taskOut_8_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_9_TREADY = task_stealSide_taskOut_9_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_10_TREADY = task_stealSide_taskOut_10_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_11_TREADY = task_stealSide_taskOut_11_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_12_TREADY = task_stealSide_taskOut_12_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_13_TREADY = task_stealSide_taskOut_13_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_14_TREADY = task_stealSide_taskOut_14_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_15_TREADY = task_stealSide_taskOut_15_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_16_TREADY = task_stealSide_taskOut_16_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_17_TREADY = task_stealSide_taskOut_17_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_18_TREADY = task_stealSide_taskOut_18_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_19_TREADY = task_stealSide_taskOut_19_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_20_TREADY = task_stealSide_taskOut_20_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_21_TREADY = task_stealSide_taskOut_21_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_22_TREADY = task_stealSide_taskOut_22_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_23_TREADY = task_stealSide_taskOut_23_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_24_TREADY = task_stealSide_taskOut_24_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_25_TREADY = task_stealSide_taskOut_25_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_26_TREADY = task_stealSide_taskOut_26_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_27_TREADY = task_stealSide_taskOut_27_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_28_TREADY = task_stealSide_taskOut_28_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_29_TREADY = task_stealSide_taskOut_29_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_30_TREADY = task_stealSide_taskOut_30_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_31_TREADY = task_stealSide_taskOut_31_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_32_TREADY = task_stealSide_taskOut_32_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_33_TREADY = task_stealSide_taskOut_33_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_34_TREADY = task_stealSide_taskOut_34_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_35_TREADY = task_stealSide_taskOut_35_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_36_TREADY = task_stealSide_taskOut_36_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_37_TREADY = task_stealSide_taskOut_37_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_38_TREADY = task_stealSide_taskOut_38_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_39_TREADY = task_stealSide_taskOut_39_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_40_TREADY = task_stealSide_taskOut_40_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_41_TREADY = task_stealSide_taskOut_41_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_42_TREADY = task_stealSide_taskOut_42_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_43_TREADY = task_stealSide_taskOut_43_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_44_TREADY = task_stealSide_taskOut_44_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_45_TREADY = task_stealSide_taskOut_45_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_46_TREADY = task_stealSide_taskOut_46_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_47_TREADY = task_stealSide_taskOut_47_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_48_TREADY = task_stealSide_taskOut_48_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_49_TREADY = task_stealSide_taskOut_49_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_50_TREADY = task_stealSide_taskOut_50_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_51_TREADY = task_stealSide_taskOut_51_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_52_TREADY = task_stealSide_taskOut_52_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_53_TREADY = task_stealSide_taskOut_53_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_54_TREADY = task_stealSide_taskOut_54_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_55_TREADY = task_stealSide_taskOut_55_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_56_TREADY = task_stealSide_taskOut_56_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_57_TREADY = task_stealSide_taskOut_57_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_58_TREADY = task_stealSide_taskOut_58_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_59_TREADY = task_stealSide_taskOut_59_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_60_TREADY = task_stealSide_taskOut_60_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_61_TREADY = task_stealSide_taskOut_61_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_62_TREADY = task_stealSide_taskOut_62_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskOut_63_TREADY = task_stealSide_taskOut_63_TREADY; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_0_TVALID = task_stealSide_taskIn_0_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_0_TDATA = task_stealSide_taskIn_0_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_1_TVALID = task_stealSide_taskIn_1_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_1_TDATA = task_stealSide_taskIn_1_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_2_TVALID = task_stealSide_taskIn_2_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_2_TDATA = task_stealSide_taskIn_2_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_3_TVALID = task_stealSide_taskIn_3_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_3_TDATA = task_stealSide_taskIn_3_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_4_TVALID = task_stealSide_taskIn_4_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_4_TDATA = task_stealSide_taskIn_4_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_5_TVALID = task_stealSide_taskIn_5_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_5_TDATA = task_stealSide_taskIn_5_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_6_TVALID = task_stealSide_taskIn_6_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_6_TDATA = task_stealSide_taskIn_6_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_7_TVALID = task_stealSide_taskIn_7_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_7_TDATA = task_stealSide_taskIn_7_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_8_TVALID = task_stealSide_taskIn_8_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_8_TDATA = task_stealSide_taskIn_8_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_9_TVALID = task_stealSide_taskIn_9_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_9_TDATA = task_stealSide_taskIn_9_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_10_TVALID = task_stealSide_taskIn_10_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_10_TDATA = task_stealSide_taskIn_10_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_11_TVALID = task_stealSide_taskIn_11_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_11_TDATA = task_stealSide_taskIn_11_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_12_TVALID = task_stealSide_taskIn_12_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_12_TDATA = task_stealSide_taskIn_12_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_13_TVALID = task_stealSide_taskIn_13_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_13_TDATA = task_stealSide_taskIn_13_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_14_TVALID = task_stealSide_taskIn_14_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_14_TDATA = task_stealSide_taskIn_14_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_15_TVALID = task_stealSide_taskIn_15_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_15_TDATA = task_stealSide_taskIn_15_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_16_TVALID = task_stealSide_taskIn_16_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_16_TDATA = task_stealSide_taskIn_16_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_17_TVALID = task_stealSide_taskIn_17_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_17_TDATA = task_stealSide_taskIn_17_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_18_TVALID = task_stealSide_taskIn_18_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_18_TDATA = task_stealSide_taskIn_18_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_19_TVALID = task_stealSide_taskIn_19_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_19_TDATA = task_stealSide_taskIn_19_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_20_TVALID = task_stealSide_taskIn_20_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_20_TDATA = task_stealSide_taskIn_20_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_21_TVALID = task_stealSide_taskIn_21_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_21_TDATA = task_stealSide_taskIn_21_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_22_TVALID = task_stealSide_taskIn_22_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_22_TDATA = task_stealSide_taskIn_22_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_23_TVALID = task_stealSide_taskIn_23_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_23_TDATA = task_stealSide_taskIn_23_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_24_TVALID = task_stealSide_taskIn_24_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_24_TDATA = task_stealSide_taskIn_24_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_25_TVALID = task_stealSide_taskIn_25_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_25_TDATA = task_stealSide_taskIn_25_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_26_TVALID = task_stealSide_taskIn_26_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_26_TDATA = task_stealSide_taskIn_26_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_27_TVALID = task_stealSide_taskIn_27_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_27_TDATA = task_stealSide_taskIn_27_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_28_TVALID = task_stealSide_taskIn_28_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_28_TDATA = task_stealSide_taskIn_28_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_29_TVALID = task_stealSide_taskIn_29_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_29_TDATA = task_stealSide_taskIn_29_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_30_TVALID = task_stealSide_taskIn_30_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_30_TDATA = task_stealSide_taskIn_30_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_31_TVALID = task_stealSide_taskIn_31_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_31_TDATA = task_stealSide_taskIn_31_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_32_TVALID = task_stealSide_taskIn_32_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_32_TDATA = task_stealSide_taskIn_32_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_33_TVALID = task_stealSide_taskIn_33_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_33_TDATA = task_stealSide_taskIn_33_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_34_TVALID = task_stealSide_taskIn_34_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_34_TDATA = task_stealSide_taskIn_34_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_35_TVALID = task_stealSide_taskIn_35_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_35_TDATA = task_stealSide_taskIn_35_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_36_TVALID = task_stealSide_taskIn_36_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_36_TDATA = task_stealSide_taskIn_36_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_37_TVALID = task_stealSide_taskIn_37_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_37_TDATA = task_stealSide_taskIn_37_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_38_TVALID = task_stealSide_taskIn_38_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_38_TDATA = task_stealSide_taskIn_38_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_39_TVALID = task_stealSide_taskIn_39_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_39_TDATA = task_stealSide_taskIn_39_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_40_TVALID = task_stealSide_taskIn_40_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_40_TDATA = task_stealSide_taskIn_40_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_41_TVALID = task_stealSide_taskIn_41_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_41_TDATA = task_stealSide_taskIn_41_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_42_TVALID = task_stealSide_taskIn_42_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_42_TDATA = task_stealSide_taskIn_42_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_43_TVALID = task_stealSide_taskIn_43_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_43_TDATA = task_stealSide_taskIn_43_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_44_TVALID = task_stealSide_taskIn_44_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_44_TDATA = task_stealSide_taskIn_44_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_45_TVALID = task_stealSide_taskIn_45_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_45_TDATA = task_stealSide_taskIn_45_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_46_TVALID = task_stealSide_taskIn_46_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_46_TDATA = task_stealSide_taskIn_46_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_47_TVALID = task_stealSide_taskIn_47_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_47_TDATA = task_stealSide_taskIn_47_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_48_TVALID = task_stealSide_taskIn_48_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_48_TDATA = task_stealSide_taskIn_48_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_49_TVALID = task_stealSide_taskIn_49_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_49_TDATA = task_stealSide_taskIn_49_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_50_TVALID = task_stealSide_taskIn_50_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_50_TDATA = task_stealSide_taskIn_50_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_51_TVALID = task_stealSide_taskIn_51_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_51_TDATA = task_stealSide_taskIn_51_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_52_TVALID = task_stealSide_taskIn_52_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_52_TDATA = task_stealSide_taskIn_52_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_53_TVALID = task_stealSide_taskIn_53_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_53_TDATA = task_stealSide_taskIn_53_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_54_TVALID = task_stealSide_taskIn_54_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_54_TDATA = task_stealSide_taskIn_54_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_55_TVALID = task_stealSide_taskIn_55_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_55_TDATA = task_stealSide_taskIn_55_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_56_TVALID = task_stealSide_taskIn_56_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_56_TDATA = task_stealSide_taskIn_56_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_57_TVALID = task_stealSide_taskIn_57_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_57_TDATA = task_stealSide_taskIn_57_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_58_TVALID = task_stealSide_taskIn_58_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_58_TDATA = task_stealSide_taskIn_58_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_59_TVALID = task_stealSide_taskIn_59_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_59_TDATA = task_stealSide_taskIn_59_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_60_TVALID = task_stealSide_taskIn_60_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_60_TDATA = task_stealSide_taskIn_60_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_61_TVALID = task_stealSide_taskIn_61_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_61_TDATA = task_stealSide_taskIn_61_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_62_TVALID = task_stealSide_taskIn_62_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_62_TDATA = task_stealSide_taskIn_62_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_63_TVALID = task_stealSide_taskIn_63_TVALID; // @[fullSysGen.scala 246:23]
  assign stealSide_io_taskIn_63_TDATA = task_stealSide_taskIn_63_TDATA; // @[fullSysGen.scala 246:23]
  assign stealSide_connSyncSide_0_ctrl_serveStealReq_valid = syncSide_connStealNtw_0_ctrl_serveStealReq_valid; // @[fullSysGen.scala 300:39]
  assign stealSide_connSyncSide_0_data_qOutTask_valid = syncSide_connStealNtw_0_data_qOutTask_valid; // @[fullSysGen.scala 300:39]
  assign stealSide_connSyncSide_0_data_qOutTask_bits = syncSide_connStealNtw_0_data_qOutTask_bits; // @[fullSysGen.scala 300:39]
  assign stealSide_connSyncSide_1_ctrl_serveStealReq_valid = syncSide_connStealNtw_1_ctrl_serveStealReq_valid; // @[fullSysGen.scala 300:39]
  assign stealSide_connSyncSide_1_data_qOutTask_valid = syncSide_connStealNtw_1_data_qOutTask_valid; // @[fullSysGen.scala 300:39]
  assign stealSide_connSyncSide_1_data_qOutTask_bits = syncSide_connStealNtw_1_data_qOutTask_bits; // @[fullSysGen.scala 300:39]
  assign continuationAllocationSide_clock = clock;
  assign continuationAllocationSide_reset = reset;
  assign continuationAllocationSide_io_contOut_0_TREADY = task_continuationAllocationSide_contOut_0_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_1_TREADY = task_continuationAllocationSide_contOut_1_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_2_TREADY = task_continuationAllocationSide_contOut_2_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_3_TREADY = task_continuationAllocationSide_contOut_3_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_4_TREADY = task_continuationAllocationSide_contOut_4_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_5_TREADY = task_continuationAllocationSide_contOut_5_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_6_TREADY = task_continuationAllocationSide_contOut_6_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_7_TREADY = task_continuationAllocationSide_contOut_7_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_8_TREADY = task_continuationAllocationSide_contOut_8_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_9_TREADY = task_continuationAllocationSide_contOut_9_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_10_TREADY = task_continuationAllocationSide_contOut_10_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_11_TREADY = task_continuationAllocationSide_contOut_11_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_12_TREADY = task_continuationAllocationSide_contOut_12_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_13_TREADY = task_continuationAllocationSide_contOut_13_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_14_TREADY = task_continuationAllocationSide_contOut_14_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_15_TREADY = task_continuationAllocationSide_contOut_15_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_16_TREADY = task_continuationAllocationSide_contOut_16_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_17_TREADY = task_continuationAllocationSide_contOut_17_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_18_TREADY = task_continuationAllocationSide_contOut_18_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_19_TREADY = task_continuationAllocationSide_contOut_19_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_20_TREADY = task_continuationAllocationSide_contOut_20_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_21_TREADY = task_continuationAllocationSide_contOut_21_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_22_TREADY = task_continuationAllocationSide_contOut_22_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_23_TREADY = task_continuationAllocationSide_contOut_23_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_24_TREADY = task_continuationAllocationSide_contOut_24_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_25_TREADY = task_continuationAllocationSide_contOut_25_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_26_TREADY = task_continuationAllocationSide_contOut_26_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_27_TREADY = task_continuationAllocationSide_contOut_27_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_28_TREADY = task_continuationAllocationSide_contOut_28_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_29_TREADY = task_continuationAllocationSide_contOut_29_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_30_TREADY = task_continuationAllocationSide_contOut_30_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_31_TREADY = task_continuationAllocationSide_contOut_31_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_32_TREADY = task_continuationAllocationSide_contOut_32_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_33_TREADY = task_continuationAllocationSide_contOut_33_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_34_TREADY = task_continuationAllocationSide_contOut_34_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_35_TREADY = task_continuationAllocationSide_contOut_35_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_36_TREADY = task_continuationAllocationSide_contOut_36_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_37_TREADY = task_continuationAllocationSide_contOut_37_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_38_TREADY = task_continuationAllocationSide_contOut_38_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_39_TREADY = task_continuationAllocationSide_contOut_39_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_40_TREADY = task_continuationAllocationSide_contOut_40_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_41_TREADY = task_continuationAllocationSide_contOut_41_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_42_TREADY = task_continuationAllocationSide_contOut_42_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_43_TREADY = task_continuationAllocationSide_contOut_43_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_44_TREADY = task_continuationAllocationSide_contOut_44_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_45_TREADY = task_continuationAllocationSide_contOut_45_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_46_TREADY = task_continuationAllocationSide_contOut_46_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_47_TREADY = task_continuationAllocationSide_contOut_47_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_48_TREADY = task_continuationAllocationSide_contOut_48_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_49_TREADY = task_continuationAllocationSide_contOut_49_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_50_TREADY = task_continuationAllocationSide_contOut_50_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_51_TREADY = task_continuationAllocationSide_contOut_51_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_52_TREADY = task_continuationAllocationSide_contOut_52_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_53_TREADY = task_continuationAllocationSide_contOut_53_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_54_TREADY = task_continuationAllocationSide_contOut_54_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_55_TREADY = task_continuationAllocationSide_contOut_55_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_56_TREADY = task_continuationAllocationSide_contOut_56_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_57_TREADY = task_continuationAllocationSide_contOut_57_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_58_TREADY = task_continuationAllocationSide_contOut_58_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_59_TREADY = task_continuationAllocationSide_contOut_59_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_60_TREADY = task_continuationAllocationSide_contOut_60_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_61_TREADY = task_continuationAllocationSide_contOut_61_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_62_TREADY = task_continuationAllocationSide_contOut_62_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_contOut_63_TREADY = task_continuationAllocationSide_contOut_63_TREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_axi_mgmt_vcas_0_ARVALID = task_continuationAllocationSide_axi_mgmt_vcas_0_ARVALID
    ; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_axi_mgmt_vcas_0_ARADDR = task_continuationAllocationSide_axi_mgmt_vcas_0_ARADDR; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_axi_mgmt_vcas_0_RREADY = task_continuationAllocationSide_axi_mgmt_vcas_0_RREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_axi_mgmt_vcas_0_AWVALID = task_continuationAllocationSide_axi_mgmt_vcas_0_AWVALID
    ; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_axi_mgmt_vcas_0_AWADDR = task_continuationAllocationSide_axi_mgmt_vcas_0_AWADDR; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_axi_mgmt_vcas_0_WVALID = task_continuationAllocationSide_axi_mgmt_vcas_0_WVALID; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_axi_mgmt_vcas_0_WDATA = task_continuationAllocationSide_axi_mgmt_vcas_0_WDATA; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_axi_mgmt_vcas_0_WSTRB = task_continuationAllocationSide_axi_mgmt_vcas_0_WSTRB; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_axi_mgmt_vcas_0_BREADY = task_continuationAllocationSide_axi_mgmt_vcas_0_BREADY; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_vcas_axi_full_0_ARREADY = task_continuationAllocationSide_vcas_axi_full_0_ARREADY
    ; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_vcas_axi_full_0_RVALID = task_continuationAllocationSide_vcas_axi_full_0_RVALID; // @[fullSysGen.scala 282:42]
  assign continuationAllocationSide_io_vcas_axi_full_0_RDATA = task_continuationAllocationSide_vcas_axi_full_0_RDATA; // @[fullSysGen.scala 282:42]
  assign syncSide_clock = clock;
  assign syncSide_reset = reset;
  assign syncSide_io_addrIn_0_TVALID = task_syncSide_addrIn_0_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_0_TDATA = task_syncSide_addrIn_0_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_1_TVALID = task_syncSide_addrIn_1_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_1_TDATA = task_syncSide_addrIn_1_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_2_TVALID = task_syncSide_addrIn_2_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_2_TDATA = task_syncSide_addrIn_2_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_3_TVALID = task_syncSide_addrIn_3_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_3_TDATA = task_syncSide_addrIn_3_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_4_TVALID = task_syncSide_addrIn_4_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_4_TDATA = task_syncSide_addrIn_4_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_5_TVALID = task_syncSide_addrIn_5_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_5_TDATA = task_syncSide_addrIn_5_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_6_TVALID = task_syncSide_addrIn_6_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_6_TDATA = task_syncSide_addrIn_6_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_7_TVALID = task_syncSide_addrIn_7_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_7_TDATA = task_syncSide_addrIn_7_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_8_TVALID = task_syncSide_addrIn_8_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_8_TDATA = task_syncSide_addrIn_8_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_9_TVALID = task_syncSide_addrIn_9_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_9_TDATA = task_syncSide_addrIn_9_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_10_TVALID = task_syncSide_addrIn_10_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_10_TDATA = task_syncSide_addrIn_10_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_11_TVALID = task_syncSide_addrIn_11_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_11_TDATA = task_syncSide_addrIn_11_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_12_TVALID = task_syncSide_addrIn_12_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_12_TDATA = task_syncSide_addrIn_12_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_13_TVALID = task_syncSide_addrIn_13_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_13_TDATA = task_syncSide_addrIn_13_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_14_TVALID = task_syncSide_addrIn_14_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_14_TDATA = task_syncSide_addrIn_14_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_15_TVALID = task_syncSide_addrIn_15_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_15_TDATA = task_syncSide_addrIn_15_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_16_TVALID = task_syncSide_addrIn_16_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_16_TDATA = task_syncSide_addrIn_16_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_17_TVALID = task_syncSide_addrIn_17_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_17_TDATA = task_syncSide_addrIn_17_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_18_TVALID = task_syncSide_addrIn_18_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_18_TDATA = task_syncSide_addrIn_18_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_19_TVALID = task_syncSide_addrIn_19_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_19_TDATA = task_syncSide_addrIn_19_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_20_TVALID = task_syncSide_addrIn_20_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_20_TDATA = task_syncSide_addrIn_20_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_21_TVALID = task_syncSide_addrIn_21_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_21_TDATA = task_syncSide_addrIn_21_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_22_TVALID = task_syncSide_addrIn_22_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_22_TDATA = task_syncSide_addrIn_22_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_23_TVALID = task_syncSide_addrIn_23_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_23_TDATA = task_syncSide_addrIn_23_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_24_TVALID = task_syncSide_addrIn_24_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_24_TDATA = task_syncSide_addrIn_24_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_25_TVALID = task_syncSide_addrIn_25_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_25_TDATA = task_syncSide_addrIn_25_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_26_TVALID = task_syncSide_addrIn_26_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_26_TDATA = task_syncSide_addrIn_26_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_27_TVALID = task_syncSide_addrIn_27_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_27_TDATA = task_syncSide_addrIn_27_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_28_TVALID = task_syncSide_addrIn_28_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_28_TDATA = task_syncSide_addrIn_28_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_29_TVALID = task_syncSide_addrIn_29_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_29_TDATA = task_syncSide_addrIn_29_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_30_TVALID = task_syncSide_addrIn_30_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_30_TDATA = task_syncSide_addrIn_30_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_31_TVALID = task_syncSide_addrIn_31_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_31_TDATA = task_syncSide_addrIn_31_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_32_TVALID = task_syncSide_addrIn_32_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_32_TDATA = task_syncSide_addrIn_32_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_33_TVALID = task_syncSide_addrIn_33_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_33_TDATA = task_syncSide_addrIn_33_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_34_TVALID = task_syncSide_addrIn_34_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_34_TDATA = task_syncSide_addrIn_34_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_35_TVALID = task_syncSide_addrIn_35_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_35_TDATA = task_syncSide_addrIn_35_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_36_TVALID = task_syncSide_addrIn_36_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_36_TDATA = task_syncSide_addrIn_36_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_37_TVALID = task_syncSide_addrIn_37_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_37_TDATA = task_syncSide_addrIn_37_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_38_TVALID = task_syncSide_addrIn_38_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_38_TDATA = task_syncSide_addrIn_38_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_39_TVALID = task_syncSide_addrIn_39_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_39_TDATA = task_syncSide_addrIn_39_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_40_TVALID = task_syncSide_addrIn_40_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_40_TDATA = task_syncSide_addrIn_40_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_41_TVALID = task_syncSide_addrIn_41_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_41_TDATA = task_syncSide_addrIn_41_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_42_TVALID = task_syncSide_addrIn_42_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_42_TDATA = task_syncSide_addrIn_42_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_43_TVALID = task_syncSide_addrIn_43_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_43_TDATA = task_syncSide_addrIn_43_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_44_TVALID = task_syncSide_addrIn_44_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_44_TDATA = task_syncSide_addrIn_44_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_45_TVALID = task_syncSide_addrIn_45_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_45_TDATA = task_syncSide_addrIn_45_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_46_TVALID = task_syncSide_addrIn_46_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_46_TDATA = task_syncSide_addrIn_46_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_47_TVALID = task_syncSide_addrIn_47_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_47_TDATA = task_syncSide_addrIn_47_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_48_TVALID = task_syncSide_addrIn_48_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_48_TDATA = task_syncSide_addrIn_48_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_49_TVALID = task_syncSide_addrIn_49_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_49_TDATA = task_syncSide_addrIn_49_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_50_TVALID = task_syncSide_addrIn_50_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_50_TDATA = task_syncSide_addrIn_50_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_51_TVALID = task_syncSide_addrIn_51_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_51_TDATA = task_syncSide_addrIn_51_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_52_TVALID = task_syncSide_addrIn_52_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_52_TDATA = task_syncSide_addrIn_52_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_53_TVALID = task_syncSide_addrIn_53_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_53_TDATA = task_syncSide_addrIn_53_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_54_TVALID = task_syncSide_addrIn_54_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_54_TDATA = task_syncSide_addrIn_54_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_55_TVALID = task_syncSide_addrIn_55_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_55_TDATA = task_syncSide_addrIn_55_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_56_TVALID = task_syncSide_addrIn_56_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_56_TDATA = task_syncSide_addrIn_56_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_57_TVALID = task_syncSide_addrIn_57_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_57_TDATA = task_syncSide_addrIn_57_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_58_TVALID = task_syncSide_addrIn_58_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_58_TDATA = task_syncSide_addrIn_58_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_59_TVALID = task_syncSide_addrIn_59_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_59_TDATA = task_syncSide_addrIn_59_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_60_TVALID = task_syncSide_addrIn_60_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_60_TDATA = task_syncSide_addrIn_60_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_61_TVALID = task_syncSide_addrIn_61_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_61_TDATA = task_syncSide_addrIn_61_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_62_TVALID = task_syncSide_addrIn_62_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_62_TDATA = task_syncSide_addrIn_62_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_63_TVALID = task_syncSide_addrIn_63_TVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_addrIn_63_TDATA = task_syncSide_addrIn_63_TDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_axi_full_argRoute_0_ARREADY = task_syncSide_axi_full_argRoute_0_ARREADY; // @[fullSysGen.scala 298:24]
  assign syncSide_io_axi_full_argRoute_0_RVALID = task_syncSide_axi_full_argRoute_0_RVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_axi_full_argRoute_0_RDATA = task_syncSide_axi_full_argRoute_0_RDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_axi_full_argRoute_0_AWREADY = task_syncSide_axi_full_argRoute_0_AWREADY; // @[fullSysGen.scala 298:24]
  assign syncSide_io_axi_full_argRoute_0_WREADY = task_syncSide_axi_full_argRoute_0_WREADY; // @[fullSysGen.scala 298:24]
  assign syncSide_io_axi_full_argRoute_0_BVALID = task_syncSide_axi_full_argRoute_0_BVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_axi_full_argRoute_1_ARREADY = task_syncSide_axi_full_argRoute_1_ARREADY; // @[fullSysGen.scala 298:24]
  assign syncSide_io_axi_full_argRoute_1_RVALID = task_syncSide_axi_full_argRoute_1_RVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_axi_full_argRoute_1_RDATA = task_syncSide_axi_full_argRoute_1_RDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_axi_full_argRoute_1_AWREADY = task_syncSide_axi_full_argRoute_1_AWREADY; // @[fullSysGen.scala 298:24]
  assign syncSide_io_axi_full_argRoute_1_WREADY = task_syncSide_axi_full_argRoute_1_WREADY; // @[fullSysGen.scala 298:24]
  assign syncSide_io_axi_full_argRoute_1_BVALID = task_syncSide_axi_full_argRoute_1_BVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_axi_full_argRoute_2_ARREADY = task_syncSide_axi_full_argRoute_2_ARREADY; // @[fullSysGen.scala 298:24]
  assign syncSide_io_axi_full_argRoute_2_RVALID = task_syncSide_axi_full_argRoute_2_RVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_axi_full_argRoute_2_RDATA = task_syncSide_axi_full_argRoute_2_RDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_io_axi_full_argRoute_3_ARREADY = task_syncSide_axi_full_argRoute_3_ARREADY; // @[fullSysGen.scala 298:24]
  assign syncSide_io_axi_full_argRoute_3_RVALID = task_syncSide_axi_full_argRoute_3_RVALID; // @[fullSysGen.scala 298:24]
  assign syncSide_io_axi_full_argRoute_3_RDATA = task_syncSide_axi_full_argRoute_3_RDATA; // @[fullSysGen.scala 298:24]
  assign syncSide_connStealNtw_0_ctrl_serveStealReq_ready = stealSide_connSyncSide_0_ctrl_serveStealReq_ready; // @[fullSysGen.scala 300:39]
  assign syncSide_connStealNtw_0_data_qOutTask_ready = stealSide_connSyncSide_0_data_qOutTask_ready; // @[fullSysGen.scala 300:39]
  assign syncSide_connStealNtw_1_ctrl_serveStealReq_ready = stealSide_connSyncSide_1_ctrl_serveStealReq_ready; // @[fullSysGen.scala 300:39]
  assign syncSide_connStealNtw_1_data_qOutTask_ready = stealSide_connSyncSide_1_data_qOutTask_ready; // @[fullSysGen.scala 300:39]
endmodule
